-- generated with romgen v3.0 by MikeJ
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity mainrom is
	port (
		clk		: in    std_logic;
		addr		: in    std_logic_vector(14 downto 0);
		data		: out   std_logic_vector(7 downto 0)
	);
end;

architecture rtl of mainrom is

	type ROM_ARRAY is array(0 to 32767) of std_logic_vector(7 downto 0);
	constant ROM : ROM_ARRAY := (
		x"F3",x"C3",x"D7",x"02",x"BF",x"1B",x"98",x"98", -- 0x0000
		x"C3",x"83",x"26",x"00",x"C3",x"B6",x"01",x"00", -- 0x0008
		x"C3",x"86",x"26",x"00",x"C3",x"D1",x"01",x"00", -- 0x0010
		x"C3",x"45",x"1B",x"00",x"C3",x"17",x"02",x"00", -- 0x0018
		x"C3",x"6A",x"14",x"00",x"C3",x"5E",x"02",x"00", -- 0x0020
		x"C3",x"89",x"26",x"11",x"11",x"00",x"00",x"00", -- 0x0028
		x"C3",x"05",x"02",x"00",x"00",x"00",x"00",x"00", -- 0x0030
		x"C3",x"3C",x"0C",x"C3",x"9D",x"04",x"C3",x"9D", -- 0x0038
		x"13",x"C3",x"77",x"05",x"C3",x"70",x"05",x"C3", -- 0x0040
		x"7F",x"05",x"C3",x"D7",x"07",x"C3",x"CD",x"07", -- 0x0048
		x"C3",x"EC",x"07",x"C3",x"DF",x"07",x"C3",x"15", -- 0x0050
		x"08",x"C3",x"0F",x"07",x"C3",x"44",x"07",x"C3", -- 0x0058
		x"4F",x"08",x"C3",x"F7",x"07",x"00",x"C3",x"98", -- 0x0060
		x"13",x"C3",x"A8",x"06",x"C3",x"0E",x"05",x"C3", -- 0x0068
		x"38",x"05",x"C3",x"D2",x"05",x"C3",x"1F",x"06", -- 0x0070
		x"C3",x"94",x"05",x"C3",x"B4",x"05",x"C3",x"02", -- 0x0078
		x"06",x"C3",x"59",x"06",x"C3",x"E4",x"06",x"C3", -- 0x0080
		x"F9",x"06",x"C3",x"04",x"07",x"C3",x"10",x"15", -- 0x0088
		x"C3",x"BD",x"04",x"C3",x"02",x"11",x"C3",x"0E", -- 0x0090
		x"11",x"C3",x"C4",x"11",x"C3",x"6A",x"0D",x"C3", -- 0x0098
		x"CB",x"10",x"C3",x"BC",x"08",x"C3",x"5D",x"08", -- 0x00A0
		x"C3",x"84",x"08",x"C3",x"9D",x"08",x"C3",x"BF", -- 0x00A8
		x"23",x"C3",x"D5",x"23",x"C3",x"CC",x"23",x"C3", -- 0x00B0
		x"6F",x"04",x"C3",x"FB",x"03",x"C3",x"F9",x"10", -- 0x00B8
		x"C3",x"13",x"11",x"C3",x"48",x"08",x"C3",x"8E", -- 0x00C0
		x"08",x"C3",x"26",x"0B",x"C3",x"15",x"0B",x"C3", -- 0x00C8
		x"2B",x"0B",x"C3",x"3B",x"08",x"C3",x"EE",x"11", -- 0x00D0
		x"C3",x"53",x"12",x"C3",x"AC",x"12",x"C3",x"73", -- 0x00D8
		x"12",x"C3",x"63",x"1A",x"C3",x"BC",x"1A",x"C3", -- 0x00E0
		x"E9",x"19",x"C3",x"F1",x"19",x"C3",x"19",x"1A", -- 0x00E8
		x"C3",x"DD",x"19",x"C3",x"84",x"13",x"C3",x"EB", -- 0x00F0
		x"14",x"C3",x"92",x"14",x"C3",x"C5",x"16",x"C3", -- 0x00F8
		x"EE",x"16",x"C3",x"5D",x"17",x"C3",x"3C",x"17", -- 0x0100
		x"C3",x"2A",x"17",x"C3",x"0A",x"17",x"C3",x"99", -- 0x0108
		x"15",x"C3",x"DF",x"15",x"C3",x"39",x"16",x"C3", -- 0x0110
		x"40",x"16",x"C3",x"76",x"16",x"C3",x"47",x"16", -- 0x0118
		x"C3",x"7E",x"16",x"C3",x"09",x"18",x"C3",x"C7", -- 0x0120
		x"18",x"C3",x"CF",x"18",x"C3",x"E4",x"18",x"C3", -- 0x0128
		x"7A",x"19",x"C3",x"3D",x"0F",x"C3",x"7A",x"0F", -- 0x0130
		x"C3",x"4C",x"14",x"C3",x"4F",x"14",x"C3",x"49", -- 0x0138
		x"14",x"C3",x"52",x"14",x"C3",x"8A",x"14",x"C3", -- 0x0140
		x"8E",x"14",x"C3",x"5F",x"14",x"C3",x"63",x"1B", -- 0x0148
		x"C3",x"70",x"14",x"C3",x"74",x"14",x"C3",x"68", -- 0x0150
		x"04",x"C3",x"FF",x"01",x"00",x"00",x"00",x"00", -- 0x0158
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0160
		x"00",x"00",x"00",x"00",x"00",x"00",x"C9",x"CD", -- 0x0168
		x"AD",x"01",x"20",x"52",x"E5",x"CD",x"99",x"01", -- 0x0170
		x"E3",x"CD",x"BE",x"7F",x"18",x"0F",x"CD",x"AD", -- 0x0178
		x"01",x"C2",x"E1",x"01",x"D1",x"E5",x"CD",x"99", -- 0x0180
		x"01",x"E3",x"CD",x"C4",x"7F",x"E3",x"F5",x"7D", -- 0x0188
		x"D3",x"A8",x"7C",x"32",x"FF",x"FF",x"F1",x"E1", -- 0x0190
		x"C9",x"F5",x"3A",x"FF",x"FF",x"2F",x"67",x"E6", -- 0x0198
		x"F3",x"32",x"FF",x"FF",x"DB",x"A8",x"6F",x"E6", -- 0x01A0
		x"F3",x"D3",x"A8",x"F1",x"C9",x"14",x"15",x"C0", -- 0x01A8
		x"47",x"7B",x"FE",x"03",x"78",x"C9",x"CD",x"7E", -- 0x01B0
		x"02",x"FA",x"6F",x"01",x"DB",x"A8",x"57",x"A1", -- 0x01B8
		x"B0",x"CD",x"80",x"F3",x"7B",x"C9",x"E5",x"CD", -- 0x01C0
		x"A3",x"02",x"E3",x"C5",x"CD",x"B6",x"01",x"18", -- 0x01C8
		x"1B",x"D5",x"CD",x"7E",x"02",x"FA",x"7E",x"01", -- 0x01D0
		x"D1",x"DB",x"A8",x"57",x"A1",x"B0",x"C3",x"85", -- 0x01D8
		x"F3",x"E3",x"E5",x"CD",x"A3",x"02",x"D1",x"E3", -- 0x01E0
		x"C5",x"CD",x"D1",x"01",x"C1",x"E3",x"F5",x"78", -- 0x01E8
		x"E6",x"3F",x"B1",x"D3",x"A8",x"7D",x"32",x"FF", -- 0x01F0
		x"FF",x"78",x"D3",x"A8",x"F1",x"E1",x"C9",x"FD", -- 0x01F8
		x"2A",x"C0",x"FC",x"18",x"12",x"E3",x"F5",x"D5", -- 0x0200
		x"7E",x"F5",x"FD",x"E1",x"23",x"5E",x"23",x"56", -- 0x0208
		x"23",x"D5",x"DD",x"E1",x"D1",x"F1",x"E3",x"D9", -- 0x0210
		x"08",x"FD",x"E5",x"F1",x"DD",x"E5",x"E1",x"CD", -- 0x0218
		x"7E",x"02",x"FA",x"2E",x"02",x"DB",x"A8",x"F5", -- 0x0220
		x"A1",x"B0",x"D9",x"C3",x"8C",x"F3",x"CD",x"A3", -- 0x0228
		x"02",x"F5",x"FD",x"E1",x"E5",x"C5",x"4F",x"06", -- 0x0230
		x"00",x"7D",x"A4",x"B2",x"21",x"C5",x"FC",x"09", -- 0x0238
		x"77",x"E5",x"08",x"D9",x"CD",x"17",x"02",x"D9", -- 0x0240
		x"08",x"E1",x"C1",x"D1",x"78",x"E6",x"3F",x"B1", -- 0x0248
		x"F3",x"D3",x"A8",x"7B",x"32",x"FF",x"FF",x"78", -- 0x0250
		x"D3",x"A8",x"73",x"08",x"D9",x"C9",x"CD",x"7E", -- 0x0258
		x"02",x"FA",x"6B",x"02",x"DB",x"A8",x"A1",x"B0", -- 0x0260
		x"D3",x"A8",x"C9",x"E5",x"CD",x"A3",x"02",x"4F", -- 0x0268
		x"06",x"00",x"7D",x"A4",x"B2",x"21",x"C5",x"FC", -- 0x0270
		x"09",x"77",x"E1",x"79",x"18",x"E0",x"F3",x"F5", -- 0x0278
		x"7C",x"07",x"07",x"E6",x"03",x"5F",x"3E",x"C0", -- 0x0280
		x"07",x"07",x"1D",x"F2",x"88",x"02",x"5F",x"2F", -- 0x0288
		x"4F",x"F1",x"F5",x"E6",x"03",x"3C",x"47",x"3E", -- 0x0290
		x"AB",x"C6",x"55",x"10",x"FC",x"57",x"A3",x"47", -- 0x0298
		x"F1",x"A7",x"C9",x"F5",x"7A",x"E6",x"C0",x"4F", -- 0x02A0
		x"F1",x"F5",x"57",x"DB",x"A8",x"47",x"E6",x"3F", -- 0x02A8
		x"B1",x"D3",x"A8",x"7A",x"0F",x"0F",x"E6",x"03", -- 0x02B0
		x"57",x"3E",x"AB",x"C6",x"55",x"15",x"F2",x"BB", -- 0x02B8
		x"02",x"A3",x"57",x"7B",x"2F",x"67",x"3A",x"FF", -- 0x02C0
		x"FF",x"2F",x"6F",x"A4",x"B2",x"32",x"FF",x"FF", -- 0x02C8
		x"78",x"D3",x"A8",x"F1",x"E6",x"03",x"C9",x"3E", -- 0x02D0
		x"82",x"D3",x"AB",x"AF",x"D3",x"A8",x"3E",x"50", -- 0x02D8
		x"D3",x"AA",x"11",x"FF",x"FF",x"AF",x"4F",x"D3", -- 0x02E0
		x"A8",x"CB",x"21",x"06",x"00",x"21",x"FF",x"FF", -- 0x02E8
		x"36",x"F0",x"7E",x"D6",x"0F",x"20",x"0B",x"77", -- 0x02F0
		x"7E",x"3C",x"20",x"06",x"04",x"CB",x"C1",x"32", -- 0x02F8
		x"FF",x"FF",x"21",x"00",x"BF",x"7E",x"2F",x"77", -- 0x0300
		x"BE",x"2F",x"77",x"20",x"07",x"2C",x"20",x"F5", -- 0x0308
		x"25",x"FA",x"05",x"03",x"2E",x"00",x"24",x"7D", -- 0x0310
		x"93",x"7C",x"9A",x"30",x"0A",x"EB",x"3A",x"FF", -- 0x0318
		x"FF",x"2F",x"6F",x"DB",x"A8",x"67",x"F9",x"78", -- 0x0320
		x"A7",x"28",x"0A",x"3A",x"FF",x"FF",x"2F",x"C6", -- 0x0328
		x"10",x"FE",x"40",x"38",x"CA",x"DB",x"A8",x"C6", -- 0x0330
		x"50",x"30",x"AC",x"21",x"00",x"00",x"39",x"7C", -- 0x0338
		x"D3",x"A8",x"7D",x"32",x"FF",x"FF",x"79",x"07", -- 0x0340
		x"07",x"07",x"07",x"4F",x"11",x"FF",x"FF",x"DB", -- 0x0348
		x"A8",x"E6",x"3F",x"D3",x"A8",x"06",x"00",x"CB", -- 0x0350
		x"01",x"30",x"0A",x"04",x"3A",x"FF",x"FF",x"2F", -- 0x0358
		x"E6",x"3F",x"32",x"FF",x"FF",x"21",x"00",x"FE", -- 0x0360
		x"7E",x"2F",x"77",x"BE",x"2F",x"77",x"20",x"09", -- 0x0368
		x"2C",x"20",x"F5",x"25",x"7C",x"FE",x"C0",x"30", -- 0x0370
		x"EF",x"2E",x"00",x"24",x"7D",x"93",x"7C",x"9A", -- 0x0378
		x"30",x"0A",x"EB",x"3A",x"FF",x"FF",x"2F",x"6F", -- 0x0380
		x"DB",x"A8",x"67",x"F9",x"78",x"A7",x"28",x"08", -- 0x0388
		x"3A",x"FF",x"FF",x"2F",x"C6",x"40",x"30",x"CA", -- 0x0390
		x"DB",x"A8",x"C6",x"40",x"30",x"B5",x"21",x"00", -- 0x0398
		x"00",x"39",x"7C",x"D3",x"A8",x"7D",x"32",x"FF", -- 0x03A0
		x"FF",x"79",x"01",x"49",x"0C",x"11",x"81",x"F3", -- 0x03A8
		x"21",x"80",x"F3",x"36",x"00",x"ED",x"B0",x"4F", -- 0x03B0
		x"06",x"04",x"21",x"C4",x"FC",x"CB",x"19",x"9F", -- 0x03B8
		x"E6",x"80",x"77",x"2B",x"10",x"F7",x"DB",x"A8", -- 0x03C0
		x"4F",x"AF",x"D3",x"A8",x"3A",x"FF",x"FF",x"2F", -- 0x03C8
		x"6F",x"3E",x"40",x"D3",x"A8",x"3A",x"FF",x"FF", -- 0x03D0
		x"2F",x"67",x"3E",x"80",x"D3",x"A8",x"3A",x"FF", -- 0x03D8
		x"FF",x"2F",x"5F",x"3E",x"C0",x"D3",x"A8",x"3A", -- 0x03E0
		x"FF",x"FF",x"2F",x"57",x"79",x"D3",x"A8",x"22", -- 0x03E8
		x"C5",x"FC",x"EB",x"22",x"C7",x"FC",x"ED",x"56", -- 0x03F0
		x"C3",x"80",x"26",x"3A",x"B1",x"FB",x"A7",x"C0", -- 0x03F8
		x"E5",x"21",x"9B",x"FC",x"F3",x"7E",x"36",x"00", -- 0x0400
		x"E1",x"FB",x"A7",x"C8",x"FE",x"03",x"28",x"1C", -- 0x0408
		x"E5",x"D5",x"C5",x"CD",x"DA",x"09",x"21",x"9B", -- 0x0410
		x"FC",x"F3",x"7E",x"36",x"00",x"FB",x"A7",x"28", -- 0x0418
		x"F8",x"F5",x"CD",x"27",x"0A",x"F1",x"C1",x"D1", -- 0x0420
		x"E1",x"FE",x"03",x"C0",x"E5",x"CD",x"68",x"04", -- 0x0428
		x"CD",x"54",x"04",x"30",x"0A",x"21",x"6A",x"FC", -- 0x0430
		x"F3",x"CD",x"F1",x"0E",x"FB",x"E1",x"C9",x"CD", -- 0x0438
		x"3B",x"08",x"3A",x"C1",x"FC",x"26",x"40",x"CD", -- 0x0440
		x"5E",x"02",x"E1",x"AF",x"ED",x"7B",x"B1",x"F6", -- 0x0448
		x"C5",x"C3",x"E6",x"63",x"3A",x"6A",x"FC",x"0F", -- 0x0450
		x"D0",x"2A",x"6B",x"FC",x"7C",x"B5",x"C8",x"2A", -- 0x0458
		x"1C",x"F4",x"23",x"7C",x"B5",x"C8",x"37",x"C9", -- 0x0460
		x"2A",x"F8",x"F3",x"22",x"FA",x"F3",x"C9",x"DB", -- 0x0468
		x"AA",x"E6",x"F0",x"F6",x"07",x"D3",x"AA",x"DB", -- 0x0470
		x"A9",x"E6",x"10",x"C0",x"DB",x"AA",x"3D",x"D3", -- 0x0478
		x"AA",x"DB",x"A9",x"E6",x"02",x"C0",x"E5",x"2A", -- 0x0480
		x"F8",x"F3",x"22",x"FA",x"F3",x"E1",x"3A",x"E1", -- 0x0488
		x"FB",x"E6",x"EF",x"32",x"E1",x"FB",x"3E",x"0D", -- 0x0490
		x"32",x"F7",x"F3",x"37",x"C9",x"3E",x"07",x"1E", -- 0x0498
		x"80",x"CD",x"02",x"11",x"3E",x"0F",x"1E",x"CF", -- 0x04A0
		x"CD",x"02",x"11",x"3E",x"0B",x"5F",x"CD",x"02", -- 0x04A8
		x"11",x"CD",x"0C",x"11",x"E6",x"40",x"32",x"AD", -- 0x04B0
		x"FC",x"3E",x"FF",x"D3",x"90",x"E5",x"D5",x"C5", -- 0x04B8
		x"F5",x"21",x"3F",x"FB",x"06",x"71",x"AF",x"77", -- 0x04C0
		x"23",x"10",x"FC",x"11",x"75",x"F9",x"06",x"7F", -- 0x04C8
		x"21",x"80",x"00",x"E5",x"D5",x"C5",x"F5",x"CD", -- 0x04D0
		x"DA",x"14",x"F1",x"C6",x"08",x"1E",x"00",x"CD", -- 0x04D8
		x"02",x"11",x"D6",x"08",x"F5",x"2E",x"0F",x"CD", -- 0x04E0
		x"77",x"14",x"EB",x"21",x"08",x"05",x"01",x"06", -- 0x04E8
		x"00",x"ED",x"B0",x"F1",x"C1",x"E1",x"D1",x"19", -- 0x04F0
		x"EB",x"3C",x"FE",x"03",x"38",x"D5",x"3E",x"07", -- 0x04F8
		x"1E",x"B8",x"CD",x"02",x"11",x"C3",x"DA",x"08", -- 0x0500
		x"04",x"04",x"78",x"88",x"FF",x"00",x"CD",x"77", -- 0x0508
		x"05",x"AF",x"32",x"AF",x"FC",x"32",x"B0",x"FC", -- 0x0510
		x"3A",x"AE",x"F3",x"32",x"B0",x"F3",x"2A",x"B3", -- 0x0518
		x"F3",x"22",x"22",x"F9",x"2A",x"B7",x"F3",x"22", -- 0x0520
		x"24",x"F9",x"CD",x"F7",x"07",x"CD",x"7E",x"07", -- 0x0528
		x"CD",x"1E",x"07",x"CD",x"94",x"05",x"18",x"38", -- 0x0530
		x"CD",x"77",x"05",x"3E",x"01",x"32",x"AF",x"FC", -- 0x0538
		x"32",x"B0",x"FC",x"3A",x"AF",x"F3",x"32",x"B0", -- 0x0540
		x"F3",x"2A",x"BD",x"F3",x"22",x"22",x"F9",x"2A", -- 0x0548
		x"C1",x"F3",x"22",x"24",x"F9",x"2A",x"C5",x"F3", -- 0x0550
		x"22",x"26",x"F9",x"2A",x"C3",x"F3",x"22",x"28", -- 0x0558
		x"F9",x"CD",x"F7",x"07",x"CD",x"7E",x"07",x"CD", -- 0x0560
		x"1E",x"07",x"CD",x"BB",x"06",x"CD",x"B4",x"05", -- 0x0568
		x"3A",x"E0",x"F3",x"F6",x"40",x"18",x"05",x"3A", -- 0x0570
		x"E0",x"F3",x"E6",x"BF",x"47",x"0E",x"01",x"78", -- 0x0578
		x"F3",x"D3",x"99",x"79",x"F6",x"80",x"D3",x"99", -- 0x0580
		x"FB",x"E5",x"78",x"06",x"00",x"21",x"DF",x"F3", -- 0x0588
		x"09",x"77",x"E1",x"C9",x"3A",x"DF",x"F3",x"E6", -- 0x0590
		x"01",x"47",x"0E",x"00",x"CD",x"7F",x"05",x"3A", -- 0x0598
		x"E0",x"F3",x"E6",x"E7",x"F6",x"10",x"47",x"0C", -- 0x05A0
		x"CD",x"7F",x"05",x"21",x"B3",x"F3",x"11",x"00", -- 0x05A8
		x"00",x"C3",x"77",x"06",x"3A",x"DF",x"F3",x"E6", -- 0x05B0
		x"01",x"47",x"0E",x"00",x"CD",x"7F",x"05",x"3A", -- 0x05B8
		x"E0",x"F3",x"E6",x"E7",x"47",x"0C",x"CD",x"7F", -- 0x05C0
		x"05",x"21",x"BD",x"F3",x"11",x"00",x"00",x"C3", -- 0x05C8
		x"77",x"06",x"CD",x"77",x"05",x"3E",x"02",x"32", -- 0x05D0
		x"AF",x"FC",x"2A",x"CF",x"F3",x"22",x"26",x"F9", -- 0x05D8
		x"2A",x"CD",x"F3",x"22",x"28",x"F9",x"2A",x"C7", -- 0x05E0
		x"F3",x"CD",x"DF",x"07",x"AF",x"06",x"03",x"D3", -- 0x05E8
		x"98",x"3C",x"20",x"FB",x"10",x"F9",x"CD",x"A1", -- 0x05F0
		x"07",x"CD",x"BB",x"06",x"CD",x"02",x"06",x"C3", -- 0x05F8
		x"70",x"05",x"3A",x"DF",x"F3",x"F6",x"02",x"47", -- 0x0600
		x"0E",x"00",x"CD",x"7F",x"05",x"3A",x"E0",x"F3", -- 0x0608
		x"E6",x"E7",x"47",x"0C",x"CD",x"7F",x"05",x"21", -- 0x0610
		x"C7",x"F3",x"11",x"03",x"7F",x"18",x"58",x"CD", -- 0x0618
		x"77",x"05",x"3E",x"03",x"32",x"AF",x"FC",x"2A", -- 0x0620
		x"D9",x"F3",x"22",x"26",x"F9",x"2A",x"D7",x"F3", -- 0x0628
		x"22",x"28",x"F9",x"2A",x"D1",x"F3",x"CD",x"DF", -- 0x0630
		x"07",x"11",x"06",x"00",x"0E",x"04",x"7A",x"06", -- 0x0638
		x"20",x"D3",x"98",x"3C",x"10",x"FB",x"0D",x"20", -- 0x0640
		x"F5",x"57",x"1D",x"20",x"EF",x"CD",x"B9",x"07", -- 0x0648
		x"CD",x"BB",x"06",x"CD",x"59",x"06",x"C3",x"70", -- 0x0650
		x"05",x"3A",x"DF",x"F3",x"E6",x"01",x"47",x"0E", -- 0x0658
		x"00",x"CD",x"7F",x"05",x"3A",x"E0",x"F3",x"E6", -- 0x0660
		x"E7",x"F6",x"08",x"47",x"0E",x"01",x"CD",x"7F", -- 0x0668
		x"05",x"21",x"D1",x"F3",x"11",x"00",x"00",x"01", -- 0x0670
		x"02",x"06",x"CD",x"90",x"06",x"06",x"0A",x"7A", -- 0x0678
		x"CD",x"91",x"06",x"06",x"05",x"7B",x"CD",x"91", -- 0x0680
		x"06",x"06",x"09",x"CD",x"90",x"06",x"06",x"05", -- 0x0688
		x"AF",x"E5",x"F5",x"7E",x"23",x"66",x"6F",x"AF", -- 0x0690
		x"29",x"8F",x"10",x"FC",x"6F",x"F1",x"B5",x"47", -- 0x0698
		x"CD",x"7F",x"05",x"E1",x"23",x"23",x"0C",x"C9", -- 0x06A0
		x"3A",x"E0",x"F3",x"47",x"0E",x"01",x"CD",x"7F", -- 0x06A8
		x"05",x"2A",x"26",x"F9",x"01",x"00",x"08",x"AF", -- 0x06B0
		x"CD",x"15",x"08",x"3A",x"E9",x"F3",x"5F",x"2A", -- 0x06B8
		x"28",x"F9",x"01",x"00",x"20",x"3E",x"D1",x"CD", -- 0x06C0
		x"CD",x"07",x"23",x"23",x"79",x"CD",x"CD",x"07", -- 0x06C8
		x"23",x"0C",x"3A",x"E0",x"F3",x"0F",x"0F",x"30", -- 0x06D0
		x"03",x"0C",x"0C",x"0C",x"7B",x"CD",x"CD",x"07", -- 0x06D8
		x"23",x"10",x"E2",x"C9",x"6F",x"26",x"00",x"29", -- 0x06E0
		x"29",x"29",x"CD",x"04",x"07",x"FE",x"08",x"28", -- 0x06E8
		x"02",x"29",x"29",x"EB",x"2A",x"26",x"F9",x"19", -- 0x06F0
		x"C9",x"6F",x"26",x"00",x"29",x"29",x"EB",x"2A", -- 0x06F8
		x"28",x"F9",x"19",x"C9",x"3A",x"E0",x"F3",x"0F", -- 0x0700
		x"0F",x"3E",x"08",x"D0",x"3E",x"20",x"C9",x"CD", -- 0x0708
		x"EC",x"07",x"E3",x"E3",x"DB",x"98",x"12",x"13", -- 0x0710
		x"0B",x"79",x"B0",x"20",x"F7",x"C9",x"CD",x"C7", -- 0x0718
		x"FD",x"2A",x"24",x"F9",x"CD",x"DF",x"07",x"3A", -- 0x0720
		x"1F",x"F9",x"2A",x"20",x"F9",x"01",x"00",x"08", -- 0x0728
		x"F5",x"F1",x"F5",x"C5",x"F3",x"CD",x"B6",x"01", -- 0x0730
		x"FB",x"C1",x"D3",x"98",x"23",x"0B",x"79",x"B0", -- 0x0738
		x"20",x"EF",x"F1",x"C9",x"EB",x"CD",x"DF",x"07", -- 0x0740
		x"1A",x"D3",x"98",x"13",x"0B",x"79",x"B0",x"20", -- 0x0748
		x"F7",x"C9",x"26",x"00",x"6F",x"29",x"29",x"29", -- 0x0750
		x"EB",x"2A",x"20",x"F9",x"19",x"11",x"40",x"FC", -- 0x0758
		x"06",x"08",x"3A",x"1F",x"F9",x"F5",x"E5",x"D5", -- 0x0760
		x"C5",x"CD",x"B6",x"01",x"FB",x"C1",x"D1",x"E1", -- 0x0768
		x"12",x"13",x"23",x"F1",x"10",x"EF",x"C9",x"CD", -- 0x0770
		x"9F",x"0B",x"28",x"25",x"30",x"3B",x"3A",x"AF", -- 0x0778
		x"FC",x"A7",x"2A",x"22",x"F9",x"01",x"C0",x"03", -- 0x0780
		x"28",x"03",x"01",x"00",x"03",x"3E",x"20",x"CD", -- 0x0788
		x"15",x"08",x"CD",x"7F",x"0A",x"21",x"B2",x"FB", -- 0x0790
		x"06",x"18",x"70",x"23",x"10",x"FC",x"C3",x"26", -- 0x0798
		x"0B",x"CD",x"32",x"08",x"01",x"00",x"18",x"C5", -- 0x07A0
		x"2A",x"C9",x"F3",x"3A",x"EA",x"F3",x"CD",x"15", -- 0x07A8
		x"08",x"2A",x"CB",x"F3",x"C1",x"AF",x"C3",x"15", -- 0x07B0
		x"08",x"CD",x"32",x"08",x"21",x"EA",x"F3",x"7E", -- 0x07B8
		x"87",x"87",x"87",x"87",x"B6",x"2A",x"D5",x"F3", -- 0x07C0
		x"01",x"00",x"06",x"18",x"E9",x"F5",x"CD",x"DF", -- 0x07C8
		x"07",x"E3",x"E3",x"F1",x"D3",x"98",x"C9",x"CD", -- 0x07D0
		x"EC",x"07",x"E3",x"E3",x"DB",x"98",x"C9",x"7D", -- 0x07D8
		x"F3",x"D3",x"99",x"7C",x"E6",x"3F",x"F6",x"40", -- 0x07E0
		x"D3",x"99",x"FB",x"C9",x"7D",x"F3",x"D3",x"99", -- 0x07E8
		x"7C",x"E6",x"3F",x"D3",x"99",x"FB",x"C9",x"3A", -- 0x07F0
		x"AF",x"FC",x"3D",x"FA",x"24",x"08",x"F5",x"CD", -- 0x07F8
		x"32",x"08",x"F1",x"C0",x"3A",x"E9",x"F3",x"87", -- 0x0800
		x"87",x"87",x"87",x"21",x"EA",x"F3",x"B6",x"2A", -- 0x0808
		x"BF",x"F3",x"01",x"20",x"00",x"F5",x"CD",x"DF", -- 0x0810
		x"07",x"F1",x"D3",x"98",x"F5",x"0B",x"79",x"B0", -- 0x0818
		x"20",x"F7",x"F1",x"C9",x"3A",x"E9",x"F3",x"87", -- 0x0820
		x"87",x"87",x"87",x"21",x"EA",x"F3",x"B6",x"47", -- 0x0828
		x"18",x"03",x"3A",x"EB",x"F3",x"47",x"0E",x"07", -- 0x0830
		x"C3",x"7F",x"05",x"CD",x"9F",x"0B",x"D8",x"3A", -- 0x0838
		x"B0",x"FC",x"CD",x"BD",x"FD",x"C3",x"4F",x"08", -- 0x0840
		x"C0",x"E5",x"CD",x"77",x"07",x"E1",x"C9",x"3D", -- 0x0848
		x"FA",x"0E",x"05",x"CA",x"38",x"05",x"3D",x"CA", -- 0x0850
		x"D2",x"05",x"C3",x"1F",x"06",x"CD",x"B6",x"FF", -- 0x0858
		x"F5",x"CD",x"6F",x"04",x"38",x"12",x"CD",x"84", -- 0x0860
		x"08",x"28",x"F6",x"F1",x"F5",x"D3",x"91",x"AF", -- 0x0868
		x"D3",x"90",x"3D",x"D3",x"90",x"F1",x"A7",x"C9", -- 0x0870
		x"AF",x"32",x"15",x"F4",x"3E",x"0D",x"CD",x"6C", -- 0x0878
		x"08",x"F1",x"37",x"C9",x"CD",x"BB",x"FF",x"DB", -- 0x0880
		x"90",x"0F",x"0F",x"3F",x"9F",x"C9",x"3E",x"1B", -- 0x0888
		x"DF",x"3E",x"59",x"DF",x"7D",x"C6",x"1F",x"DF", -- 0x0890
		x"7C",x"C6",x"1F",x"DF",x"C9",x"E5",x"F5",x"21", -- 0x0898
		x"A6",x"FC",x"AF",x"BE",x"77",x"28",x"0D",x"F1", -- 0x08A0
		x"D6",x"40",x"FE",x"20",x"38",x"04",x"C6",x"40", -- 0x08A8
		x"BF",x"37",x"E1",x"C9",x"F1",x"FE",x"01",x"20", -- 0x08B0
		x"F7",x"77",x"E1",x"C9",x"E5",x"D5",x"C5",x"F5", -- 0x08B8
		x"CD",x"A4",x"FD",x"CD",x"9F",x"0B",x"30",x"12", -- 0x08C0
		x"CD",x"2E",x"0A",x"F1",x"F5",x"CD",x"DF",x"08", -- 0x08C8
		x"CD",x"E1",x"09",x"3A",x"DD",x"F3",x"3D",x"32", -- 0x08D0
		x"61",x"F6",x"F1",x"C1",x"D1",x"E1",x"C9",x"CD", -- 0x08D8
		x"9D",x"08",x"D0",x"4F",x"20",x"0D",x"21",x"A7", -- 0x08E0
		x"FC",x"7E",x"A7",x"C2",x"8F",x"09",x"79",x"FE", -- 0x08E8
		x"20",x"38",x"21",x"2A",x"DC",x"F3",x"FE",x"7F", -- 0x08F0
		x"CA",x"E3",x"0A",x"CD",x"E6",x"0B",x"CD",x"44", -- 0x08F8
		x"0A",x"C0",x"AF",x"CD",x"2B",x"0C",x"26",x"01", -- 0x0900
		x"CD",x"61",x"0A",x"C0",x"CD",x"69",x"0A",x"2E", -- 0x0908
		x"01",x"C3",x"88",x"0A",x"21",x"2D",x"09",x"0E", -- 0x0910
		x"0C",x"23",x"23",x"A7",x"0D",x"F8",x"BE",x"23", -- 0x0918
		x"20",x"F7",x"4E",x"23",x"46",x"2A",x"DC",x"F3", -- 0x0920
		x"CD",x"2D",x"09",x"AF",x"C9",x"C5",x"C9",x"07", -- 0x0928
		x"13",x"11",x"08",x"4C",x"0A",x"09",x"71",x"0A", -- 0x0930
		x"0A",x"08",x"09",x"0B",x"7F",x"0A",x"0C",x"7E", -- 0x0938
		x"07",x"0D",x"81",x"0A",x"1B",x"89",x"09",x"1C", -- 0x0940
		x"5B",x"0A",x"1D",x"4C",x"0A",x"1E",x"57",x"0A", -- 0x0948
		x"1F",x"61",x"0A",x"6A",x"7E",x"07",x"45",x"7E", -- 0x0950
		x"07",x"4B",x"EE",x"0A",x"4A",x"05",x"0B",x"6C", -- 0x0958
		x"EC",x"0A",x"4C",x"B4",x"0A",x"4D",x"85",x"0A", -- 0x0960
		x"59",x"86",x"09",x"41",x"57",x"0A",x"42",x"61", -- 0x0968
		x"0A",x"43",x"44",x"0A",x"44",x"55",x"0A",x"48", -- 0x0970
		x"7F",x"0A",x"78",x"80",x"09",x"79",x"83",x"09", -- 0x0978
		x"3E",x"01",x"01",x"3E",x"02",x"01",x"3E",x"04", -- 0x0980
		x"01",x"3E",x"FF",x"32",x"A7",x"FC",x"C9",x"F2", -- 0x0988
		x"9D",x"09",x"36",x"00",x"79",x"21",x"51",x"09", -- 0x0990
		x"0E",x"0F",x"C3",x"19",x"09",x"3D",x"28",x"1E", -- 0x0998
		x"3D",x"28",x"25",x"3D",x"77",x"3A",x"B0",x"F3", -- 0x09A0
		x"11",x"DD",x"F3",x"28",x"06",x"36",x"03",x"CD", -- 0x09A8
		x"32",x"0C",x"1B",x"47",x"79",x"D6",x"20",x"B8", -- 0x09B0
		x"3C",x"12",x"D8",x"78",x"12",x"C9",x"77",x"79", -- 0x09B8
		x"D6",x"34",x"28",x"0B",x"3D",x"28",x"0F",x"C9", -- 0x09C0
		x"77",x"79",x"D6",x"34",x"20",x"05",x"3C",x"32", -- 0x09C8
		x"AA",x"FC",x"C9",x"3D",x"C0",x"3C",x"32",x"A9", -- 0x09D0
		x"FC",x"C9",x"3A",x"A9",x"FC",x"A7",x"C0",x"18", -- 0x09D8
		x"05",x"3A",x"A9",x"FC",x"A7",x"C8",x"CD",x"A9", -- 0x09E0
		x"FD",x"CD",x"9F",x"0B",x"D0",x"2A",x"DC",x"F3", -- 0x09E8
		x"E5",x"CD",x"D8",x"0B",x"32",x"CC",x"FB",x"6F", -- 0x09F0
		x"26",x"00",x"29",x"29",x"29",x"EB",x"2A",x"24", -- 0x09F8
		x"F9",x"E5",x"19",x"CD",x"A5",x"0B",x"21",x"1F", -- 0x0A00
		x"FC",x"06",x"08",x"3A",x"AA",x"FC",x"A7",x"28", -- 0x0A08
		x"02",x"06",x"03",x"7E",x"2F",x"77",x"2B",x"10", -- 0x0A10
		x"FA",x"E1",x"01",x"F8",x"07",x"09",x"CD",x"BE", -- 0x0A18
		x"0B",x"E1",x"0E",x"FF",x"C3",x"E6",x"0B",x"3A", -- 0x0A20
		x"A9",x"FC",x"A7",x"C0",x"18",x"05",x"3A",x"A9", -- 0x0A28
		x"FC",x"A7",x"C8",x"CD",x"AE",x"FD",x"CD",x"9F", -- 0x0A30
		x"0B",x"D0",x"2A",x"DC",x"F3",x"3A",x"CC",x"FB", -- 0x0A38
		x"4F",x"C3",x"E6",x"0B",x"3A",x"B0",x"F3",x"BC", -- 0x0A40
		x"C8",x"24",x"18",x"1D",x"CD",x"55",x"0A",x"C0", -- 0x0A48
		x"3A",x"B0",x"F3",x"67",x"11",x"25",x"3E",x"2D", -- 0x0A50
		x"C8",x"18",x"0E",x"CD",x"44",x"0A",x"C0",x"26", -- 0x0A58
		x"01",x"CD",x"32",x"0C",x"BD",x"C8",x"38",x"05", -- 0x0A60
		x"2C",x"22",x"DC",x"F3",x"C9",x"2D",x"AF",x"18", -- 0x0A68
		x"F8",x"3E",x"20",x"CD",x"DF",x"08",x"3A",x"DD", -- 0x0A70
		x"F3",x"3D",x"E6",x"07",x"20",x"F3",x"C9",x"2E", -- 0x0A78
		x"01",x"26",x"01",x"18",x"E4",x"CD",x"81",x"0A", -- 0x0A80
		x"CD",x"32",x"0C",x"95",x"D8",x"CA",x"EC",x"0A", -- 0x0A88
		x"E5",x"F5",x"4F",x"06",x"00",x"CD",x"1D",x"0C", -- 0x0A90
		x"6B",x"62",x"23",x"ED",x"B0",x"21",x"CA",x"FB", -- 0x0A98
		x"35",x"F1",x"E1",x"F5",x"2C",x"CD",x"AA",x"0B", -- 0x0AA0
		x"2D",x"CD",x"C3",x"0B",x"2C",x"F1",x"3D",x"20", -- 0x0AA8
		x"F2",x"C3",x"EC",x"0A",x"CD",x"81",x"0A",x"CD", -- 0x0AB0
		x"32",x"0C",x"67",x"95",x"D8",x"CA",x"EC",x"0A", -- 0x0AB8
		x"6C",x"E5",x"F5",x"4F",x"06",x"00",x"CD",x"1D", -- 0x0AC0
		x"0C",x"6B",x"62",x"E5",x"2B",x"ED",x"B8",x"E1", -- 0x0AC8
		x"74",x"F1",x"E1",x"F5",x"2D",x"CD",x"AA",x"0B", -- 0x0AD0
		x"2C",x"CD",x"C3",x"0B",x"2D",x"F1",x"3D",x"20", -- 0x0AD8
		x"F2",x"18",x"09",x"CD",x"4C",x"0A",x"C8",x"0E", -- 0x0AE0
		x"20",x"C3",x"E6",x"0B",x"26",x"01",x"CD",x"29", -- 0x0AE8
		x"0C",x"E5",x"CD",x"F2",x"0B",x"CD",x"DF",x"07", -- 0x0AF0
		x"E1",x"3E",x"20",x"D3",x"98",x"24",x"3A",x"B0", -- 0x0AF8
		x"F3",x"BC",x"30",x"F5",x"C9",x"E5",x"CD",x"EE", -- 0x0B00
		x"0A",x"E1",x"CD",x"32",x"0C",x"BD",x"D8",x"C8", -- 0x0B08
		x"26",x"01",x"2C",x"18",x"F0",x"CD",x"B8",x"FD", -- 0x0B10
		x"AF",x"CD",x"9C",x"0B",x"D0",x"E5",x"2A",x"B1", -- 0x0B18
		x"F3",x"CD",x"EC",x"0A",x"E1",x"C9",x"3A",x"DE", -- 0x0B20
		x"F3",x"A7",x"C8",x"CD",x"B3",x"FD",x"3E",x"FF", -- 0x0B28
		x"CD",x"9C",x"0B",x"D0",x"E5",x"3A",x"DC",x"F3", -- 0x0B30
		x"21",x"B1",x"F3",x"BE",x"3E",x"0A",x"20",x"01", -- 0x0B38
		x"DF",x"3A",x"EB",x"FB",x"0F",x"21",x"7F",x"F8", -- 0x0B40
		x"3E",x"01",x"38",x"04",x"21",x"CF",x"F8",x"AF", -- 0x0B48
		x"32",x"CD",x"FB",x"11",x"18",x"FC",x"D5",x"06", -- 0x0B50
		x"28",x"3E",x"20",x"12",x"13",x"10",x"FC",x"D1", -- 0x0B58
		x"0E",x"05",x"3A",x"B0",x"F3",x"D6",x"04",x"38", -- 0x0B60
		x"2B",x"06",x"FF",x"04",x"D6",x"05",x"30",x"FB", -- 0x0B68
		x"78",x"A7",x"28",x"20",x"3E",x"13",x"C5",x"0E", -- 0x0B70
		x"00",x"7E",x"23",x"0C",x"CD",x"9D",x"08",x"30", -- 0x0B78
		x"F8",x"20",x"04",x"FE",x"20",x"38",x"01",x"12", -- 0x0B80
		x"13",x"10",x"EE",x"3E",x"10",x"91",x"4F",x"09", -- 0x0B88
		x"C1",x"0D",x"20",x"E1",x"2A",x"B1",x"F3",x"CD", -- 0x0B90
		x"C3",x"0B",x"E1",x"C9",x"32",x"DE",x"F3",x"3A", -- 0x0B98
		x"AF",x"FC",x"FE",x"02",x"C9",x"E5",x"0E",x"08", -- 0x0BA0
		x"18",x"0A",x"E5",x"26",x"01",x"CD",x"F2",x"0B", -- 0x0BA8
		x"3A",x"B0",x"F3",x"4F",x"06",x"00",x"11",x"18", -- 0x0BB0
		x"FC",x"CD",x"0F",x"07",x"E1",x"C9",x"E5",x"0E", -- 0x0BB8
		x"08",x"18",x"0A",x"E5",x"26",x"01",x"CD",x"F2", -- 0x0BC0
		x"0B",x"3A",x"B0",x"F3",x"4F",x"06",x"00",x"EB", -- 0x0BC8
		x"21",x"18",x"FC",x"CD",x"44",x"07",x"E1",x"C9", -- 0x0BD0
		x"E5",x"CD",x"F2",x"0B",x"CD",x"EC",x"07",x"E3", -- 0x0BD8
		x"E3",x"DB",x"98",x"4F",x"E1",x"C9",x"E5",x"CD", -- 0x0BE0
		x"F2",x"0B",x"CD",x"DF",x"07",x"79",x"D3",x"98", -- 0x0BE8
		x"E1",x"C9",x"C5",x"5C",x"26",x"00",x"54",x"2D", -- 0x0BF0
		x"29",x"29",x"29",x"4D",x"44",x"29",x"29",x"19", -- 0x0BF8
		x"3A",x"AF",x"FC",x"A7",x"3A",x"B0",x"F3",x"28", -- 0x0C00
		x"04",x"D6",x"22",x"18",x"03",x"09",x"D6",x"2A", -- 0x0C08
		x"2F",x"A7",x"1F",x"5F",x"19",x"EB",x"2A",x"22", -- 0x0C10
		x"F9",x"19",x"2B",x"C1",x"C9",x"E5",x"11",x"B1", -- 0x0C18
		x"FB",x"26",x"00",x"19",x"7E",x"EB",x"E1",x"A7", -- 0x0C20
		x"C9",x"3E",x"AF",x"F5",x"CD",x"1D",x"0C",x"F1", -- 0x0C28
		x"12",x"C9",x"3A",x"DE",x"F3",x"E5",x"21",x"B1", -- 0x0C30
		x"F3",x"86",x"E1",x"C9",x"E5",x"D5",x"C5",x"F5", -- 0x0C38
		x"D9",x"08",x"E5",x"D5",x"C5",x"F5",x"FD",x"E5", -- 0x0C40
		x"DD",x"E5",x"CD",x"9A",x"FD",x"DB",x"99",x"A7", -- 0x0C48
		x"F2",x"02",x"0D",x"CD",x"9F",x"FD",x"FB",x"32", -- 0x0C50
		x"E7",x"F3",x"E6",x"20",x"21",x"6D",x"FC",x"C4", -- 0x0C58
		x"F1",x"0E",x"2A",x"A2",x"FC",x"2B",x"7C",x"B5", -- 0x0C60
		x"20",x"09",x"21",x"7F",x"FC",x"CD",x"F1",x"0E", -- 0x0C68
		x"2A",x"A0",x"FC",x"22",x"A2",x"FC",x"2A",x"9E", -- 0x0C70
		x"FC",x"23",x"22",x"9E",x"FC",x"3A",x"3F",x"FB", -- 0x0C78
		x"4F",x"AF",x"CB",x"19",x"F5",x"C5",x"DC",x"3B", -- 0x0C80
		x"11",x"C1",x"F1",x"3C",x"FE",x"03",x"38",x"F2", -- 0x0C88
		x"21",x"F6",x"F3",x"35",x"20",x"6C",x"36",x"03", -- 0x0C90
		x"AF",x"CD",x"0C",x"12",x"E6",x"30",x"F5",x"3E", -- 0x0C98
		x"01",x"CD",x"0C",x"12",x"E6",x"30",x"07",x"07", -- 0x0CA0
		x"C1",x"B0",x"F5",x"CD",x"26",x"12",x"E6",x"01", -- 0x0CA8
		x"C1",x"B0",x"4F",x"21",x"E8",x"F3",x"AE",x"A6", -- 0x0CB0
		x"71",x"4F",x"0F",x"21",x"70",x"FC",x"DC",x"F1", -- 0x0CB8
		x"0E",x"CB",x"11",x"21",x"7C",x"FC",x"DC",x"F1", -- 0x0CC0
		x"0E",x"CB",x"11",x"21",x"76",x"FC",x"DC",x"F1", -- 0x0CC8
		x"0E",x"CB",x"11",x"21",x"79",x"FC",x"DC",x"F1", -- 0x0CD0
		x"0E",x"CB",x"11",x"21",x"73",x"FC",x"DC",x"F1", -- 0x0CD8
		x"0E",x"AF",x"32",x"D9",x"FB",x"CD",x"12",x"0D", -- 0x0CE0
		x"20",x"18",x"21",x"F7",x"F3",x"35",x"20",x"12", -- 0x0CE8
		x"36",x"01",x"21",x"DA",x"FB",x"11",x"DB",x"FB", -- 0x0CF0
		x"01",x"0A",x"00",x"36",x"FF",x"ED",x"B0",x"CD", -- 0x0CF8
		x"4E",x"0D",x"DD",x"E1",x"FD",x"E1",x"F1",x"C1", -- 0x0D00
		x"D1",x"E1",x"08",x"D9",x"F1",x"C1",x"D1",x"E1", -- 0x0D08
		x"FB",x"C9",x"DB",x"AA",x"E6",x"F0",x"4F",x"06", -- 0x0D10
		x"0B",x"21",x"E5",x"FB",x"79",x"D3",x"AA",x"DB", -- 0x0D18
		x"A9",x"77",x"0C",x"23",x"10",x"F6",x"3A",x"B0", -- 0x0D20
		x"FB",x"A7",x"28",x"0E",x"3A",x"EB",x"FB",x"FE", -- 0x0D28
		x"E8",x"20",x"07",x"DD",x"21",x"9B",x"40",x"C3", -- 0x0D30
		x"FF",x"01",x"11",x"E5",x"FB",x"06",x"0B",x"1B", -- 0x0D38
		x"2B",x"1A",x"BE",x"20",x"04",x"10",x"F8",x"18", -- 0x0D40
		x"05",x"3E",x"0D",x"32",x"F7",x"F3",x"06",x"0B", -- 0x0D48
		x"21",x"DA",x"FB",x"11",x"E5",x"FB",x"1A",x"4F", -- 0x0D50
		x"AE",x"A6",x"71",x"C4",x"89",x"0D",x"13",x"23", -- 0x0D58
		x"10",x"F4",x"2A",x"FA",x"F3",x"3A",x"F8",x"F3", -- 0x0D60
		x"95",x"C9",x"FB",x"E5",x"D5",x"C5",x"CD",x"9F", -- 0x0D68
		x"0B",x"30",x"0F",x"3A",x"CD",x"FB",x"21",x"EB", -- 0x0D70
		x"FB",x"AE",x"21",x"DE",x"F3",x"A6",x"0F",x"DC", -- 0x0D78
		x"2B",x"0B",x"CD",x"62",x"0D",x"C1",x"D1",x"E1", -- 0x0D80
		x"C9",x"E5",x"D5",x"C5",x"F5",x"3E",x"0B",x"90", -- 0x0D88
		x"87",x"87",x"87",x"4F",x"06",x"08",x"F1",x"1F", -- 0x0D90
		x"C5",x"F5",x"DC",x"21",x"10",x"F1",x"C1",x"0C", -- 0x0D98
		x"10",x"F5",x"C3",x"DB",x"08",x"30",x"31",x"32", -- 0x0DA0
		x"33",x"34",x"35",x"36",x"37",x"38",x"39",x"2D", -- 0x0DA8
		x"3D",x"5C",x"5B",x"5D",x"3B",x"27",x"60",x"2C", -- 0x0DB0
		x"2E",x"2F",x"FF",x"61",x"62",x"63",x"64",x"65", -- 0x0DB8
		x"66",x"67",x"68",x"69",x"6A",x"6B",x"6C",x"6D", -- 0x0DC0
		x"6E",x"6F",x"70",x"71",x"72",x"73",x"74",x"75", -- 0x0DC8
		x"76",x"77",x"78",x"79",x"7A",x"29",x"21",x"40", -- 0x0DD0
		x"23",x"24",x"25",x"5E",x"26",x"2A",x"28",x"5F", -- 0x0DD8
		x"2B",x"7C",x"7B",x"7D",x"3A",x"22",x"7E",x"3C", -- 0x0DE0
		x"3E",x"3F",x"FF",x"41",x"42",x"43",x"44",x"45", -- 0x0DE8
		x"46",x"47",x"48",x"49",x"4A",x"4B",x"4C",x"4D", -- 0x0DF0
		x"4E",x"4F",x"50",x"51",x"52",x"53",x"54",x"55", -- 0x0DF8
		x"56",x"57",x"58",x"59",x"5A",x"09",x"AC",x"AB", -- 0x0E00
		x"BA",x"EF",x"BD",x"F4",x"FB",x"EC",x"07",x"17", -- 0x0E08
		x"F1",x"1E",x"01",x"0D",x"06",x"05",x"BB",x"F3", -- 0x0E10
		x"F2",x"1D",x"FF",x"C4",x"11",x"BC",x"C7",x"CD", -- 0x0E18
		x"14",x"15",x"13",x"DC",x"C6",x"DD",x"C8",x"0B", -- 0x0E20
		x"1B",x"C2",x"DB",x"CC",x"18",x"D2",x"12",x"C0", -- 0x0E28
		x"1A",x"CF",x"1C",x"19",x"0F",x"0A",x"00",x"FD", -- 0x0E30
		x"FC",x"00",x"00",x"F5",x"00",x"00",x"08",x"1F", -- 0x0E38
		x"F0",x"16",x"02",x"0E",x"04",x"03",x"F7",x"AE", -- 0x0E40
		x"AF",x"F6",x"FF",x"FE",x"00",x"FA",x"C1",x"CE", -- 0x0E48
		x"D4",x"10",x"D6",x"DF",x"CA",x"DE",x"C9",x"0C", -- 0x0E50
		x"D3",x"C3",x"D7",x"CB",x"A9",x"D1",x"00",x"C5", -- 0x0E58
		x"D5",x"D0",x"F9",x"AA",x"F8",x"EB",x"9F",x"D9", -- 0x0E60
		x"BF",x"9B",x"98",x"E0",x"E1",x"E7",x"87",x"EE", -- 0x0E68
		x"E9",x"00",x"ED",x"DA",x"B7",x"B9",x"E5",x"86", -- 0x0E70
		x"A6",x"A7",x"FF",x"84",x"97",x"8D",x"8B",x"8C", -- 0x0E78
		x"94",x"81",x"B1",x"A1",x"91",x"B3",x"B5",x"E6", -- 0x0E80
		x"A4",x"A2",x"A3",x"83",x"93",x"89",x"96",x"82", -- 0x0E88
		x"95",x"88",x"8A",x"A0",x"85",x"D8",x"AD",x"9E", -- 0x0E90
		x"BE",x"9C",x"9D",x"00",x"00",x"E2",x"80",x"00", -- 0x0E98
		x"00",x"00",x"E8",x"EA",x"B6",x"B8",x"E4",x"8F", -- 0x0EA0
		x"00",x"A8",x"FF",x"8E",x"00",x"00",x"00",x"00", -- 0x0EA8
		x"99",x"9A",x"B0",x"00",x"92",x"B2",x"B4",x"00", -- 0x0EB0
		x"A5",x"00",x"E3",x"00",x"00",x"00",x"00",x"90", -- 0x0EB8
		x"00",x"00",x"00",x"00",x"00",x"59",x"16",x"00", -- 0x0EC0
		x"21",x"99",x"FB",x"19",x"7E",x"A7",x"20",x"13", -- 0x0EC8
		x"EB",x"29",x"29",x"29",x"29",x"11",x"2F",x"F5", -- 0x0ED0
		x"19",x"EB",x"1A",x"A7",x"C8",x"CD",x"55",x"0F", -- 0x0ED8
		x"13",x"18",x"F7",x"2A",x"1C",x"F4",x"23",x"7C", -- 0x0EE0
		x"B5",x"28",x"E5",x"21",x"AD",x"FB",x"19",x"19", -- 0x0EE8
		x"19",x"7E",x"E6",x"01",x"C8",x"7E",x"F6",x"04", -- 0x0EF0
		x"BE",x"C8",x"77",x"EE",x"05",x"C0",x"3A",x"D8", -- 0x0EF8
		x"FB",x"3C",x"32",x"D8",x"FB",x"C9",x"3A",x"EB", -- 0x0F00
		x"FB",x"0F",x"3E",x"0C",x"DE",x"00",x"18",x"45", -- 0x0F08
		x"CD",x"D1",x"FD",x"5F",x"16",x"00",x"21",x"03", -- 0x0F10
		x"10",x"19",x"7E",x"A7",x"C8",x"18",x"36",x"3A", -- 0x0F18
		x"EB",x"FB",x"5F",x"F6",x"FE",x"CB",x"63",x"20", -- 0x0F20
		x"02",x"E6",x"FD",x"2F",x"3C",x"32",x"AC",x"FC", -- 0x0F28
		x"18",x"32",x"00",x"00",x"00",x"00",x"21",x"AB", -- 0x0F30
		x"FC",x"7E",x"2F",x"77",x"2F",x"A7",x"3E",x"0C", -- 0x0F38
		x"28",x"01",x"3C",x"D3",x"AB",x"C9",x"3A",x"EB", -- 0x0F40
		x"FB",x"0F",x"0F",x"3E",x"03",x"30",x"01",x"3C", -- 0x0F48
		x"32",x"9B",x"FC",x"38",x"0F",x"2A",x"F8",x"F3", -- 0x0F50
		x"77",x"CD",x"5B",x"10",x"3A",x"FA",x"F3",x"BD", -- 0x0F58
		x"C8",x"22",x"F8",x"F3",x"3A",x"DB",x"F3",x"A7", -- 0x0F60
		x"C8",x"3A",x"D9",x"FB",x"A7",x"C0",x"3E",x"0F", -- 0x0F68
		x"32",x"D9",x"FB",x"D3",x"AB",x"3E",x"0A",x"3D", -- 0x0F70
		x"20",x"FD",x"A7",x"3E",x"0E",x"28",x"01",x"3C", -- 0x0F78
		x"D3",x"AB",x"C9",x"3A",x"EB",x"FB",x"5F",x"1F", -- 0x0F80
		x"1F",x"F5",x"7B",x"2F",x"30",x"10",x"1F",x"1F", -- 0x0F88
		x"07",x"E6",x"03",x"CB",x"4F",x"20",x"09",x"CB", -- 0x0F90
		x"63",x"20",x"05",x"F6",x"04",x"11",x"E6",x"01", -- 0x0F98
		x"5F",x"87",x"83",x"87",x"87",x"87",x"87",x"5F", -- 0x0FA0
		x"16",x"00",x"21",x"A5",x"0D",x"19",x"42",x"09", -- 0x0FA8
		x"F1",x"7E",x"3C",x"CA",x"1F",x"0F",x"3D",x"C8", -- 0x0FB0
		x"38",x"16",x"E6",x"DF",x"D6",x"40",x"FE",x"20", -- 0x0FB8
		x"D0",x"18",x"92",x"3A",x"EB",x"FB",x"0F",x"38", -- 0x0FC0
		x"04",x"79",x"C6",x"05",x"4F",x"C3",x"C5",x"0E", -- 0x0FC8
		x"FE",x"20",x"30",x"0B",x"F5",x"3E",x"01",x"CD", -- 0x0FD0
		x"55",x"0F",x"F1",x"C6",x"40",x"18",x"E2",x"21", -- 0x0FD8
		x"AB",x"FC",x"34",x"35",x"28",x"0A",x"FE",x"61", -- 0x0FE0
		x"38",x"27",x"FE",x"7B",x"30",x"23",x"E6",x"DF", -- 0x0FE8
		x"ED",x"5B",x"AC",x"FC",x"1C",x"1D",x"28",x"C9", -- 0x0FF0
		x"57",x"F6",x"20",x"21",x"66",x"10",x"0E",x"06", -- 0x0FF8
		x"ED",x"B9",x"7A",x"20",x"BC",x"23",x"0E",x"06", -- 0x1000
		x"09",x"1D",x"20",x"FC",x"7E",x"CB",x"6A",x"20", -- 0x1008
		x"B0",x"0E",x"1F",x"21",x"9D",x"10",x"ED",x"B9", -- 0x1010
		x"20",x"A7",x"0E",x"1F",x"23",x"09",x"7E",x"18", -- 0x1018
		x"A0",x"79",x"21",x"96",x"1B",x"CD",x"CC",x"FD", -- 0x1020
		x"16",x"0F",x"BE",x"23",x"5E",x"23",x"D5",x"D8", -- 0x1028
		x"D1",x"18",x"F7",x"00",x"00",x"00",x"00",x"00", -- 0x1030
		x"00",x"00",x"00",x"00",x"00",x"1B",x"09",x"00", -- 0x1038
		x"08",x"18",x"0D",x"20",x"0C",x"12",x"7F",x"1D", -- 0x1040
		x"1E",x"1F",x"1C",x"2A",x"2B",x"2F",x"30",x"31", -- 0x1048
		x"32",x"33",x"34",x"35",x"36",x"37",x"38",x"39", -- 0x1050
		x"2D",x"2C",x"2E",x"AF",x"32",x"AC",x"FC",x"18", -- 0x1058
		x"61",x"61",x"65",x"69",x"6F",x"75",x"79",x"85", -- 0x1060
		x"8A",x"8D",x"95",x"97",x"79",x"A0",x"82",x"A1", -- 0x1068
		x"A2",x"A3",x"79",x"83",x"88",x"8C",x"93",x"96", -- 0x1070
		x"79",x"84",x"89",x"8B",x"94",x"81",x"98",x"83", -- 0x1078
		x"88",x"8C",x"93",x"96",x"84",x"89",x"8B",x"94", -- 0x1080
		x"81",x"98",x"A0",x"82",x"A1",x"A2",x"A3",x"85", -- 0x1088
		x"8A",x"8D",x"95",x"97",x"B1",x"B3",x"B5",x"B7", -- 0x1090
		x"A4",x"86",x"87",x"91",x"B9",x"79",x"41",x"45", -- 0x1098
		x"49",x"4F",x"55",x"8E",x"45",x"49",x"99",x"9A", -- 0x10A0
		x"59",x"41",x"90",x"49",x"4F",x"55",x"41",x"45", -- 0x10A8
		x"49",x"4F",x"55",x"B0",x"B2",x"B4",x"B6",x"A5", -- 0x10B0
		x"8F",x"80",x"92",x"B8",x"59",x"00",x"00",x"00", -- 0x10B8
		x"00",x"00",x"23",x"7D",x"FE",x"18",x"C0",x"21", -- 0x10C0
		x"F0",x"FB",x"C9",x"E5",x"D5",x"C5",x"CD",x"C2", -- 0x10C8
		x"FD",x"CD",x"6A",x"0D",x"20",x"0B",x"CD",x"DA", -- 0x10D0
		x"09",x"CD",x"6A",x"0D",x"28",x"FB",x"CD",x"27", -- 0x10D8
		x"0A",x"21",x"9B",x"FC",x"7E",x"FE",x"04",x"20", -- 0x10E0
		x"02",x"36",x"00",x"2A",x"FA",x"F3",x"4E",x"CD", -- 0x10E8
		x"C2",x"10",x"22",x"FA",x"F3",x"79",x"C3",x"DB", -- 0x10F0
		x"08",x"E5",x"21",x"00",x"00",x"CD",x"FB",x"03", -- 0x10F8
		x"E1",x"C9",x"F3",x"D3",x"A0",x"F5",x"7B",x"D3", -- 0x1100
		x"A1",x"FB",x"F1",x"C9",x"3E",x"0E",x"D3",x"A0", -- 0x1108
		x"DB",x"A2",x"C9",x"AF",x"1E",x"55",x"CD",x"02", -- 0x1110
		x"11",x"5F",x"3C",x"CD",x"02",x"11",x"1E",x"BE", -- 0x1118
		x"3E",x"07",x"CD",x"02",x"11",x"5F",x"3C",x"CD", -- 0x1120
		x"02",x"11",x"01",x"D0",x"07",x"CD",x"33",x"11", -- 0x1128
		x"C3",x"BD",x"04",x"0B",x"E3",x"E3",x"78",x"B1", -- 0x1130
		x"20",x"F9",x"C9",x"47",x"CD",x"70",x"14",x"2B", -- 0x1138
		x"56",x"2B",x"5E",x"1B",x"73",x"23",x"72",x"7A", -- 0x1140
		x"B3",x"C0",x"78",x"32",x"3E",x"FB",x"CD",x"E2", -- 0x1148
		x"11",x"FE",x"FF",x"28",x"5B",x"57",x"E6",x"E0", -- 0x1150
		x"07",x"07",x"07",x"4F",x"7A",x"E6",x"1F",x"77", -- 0x1158
		x"CD",x"E2",x"11",x"2B",x"77",x"0C",x"0D",x"C8", -- 0x1160
		x"CD",x"E2",x"11",x"57",x"E6",x"C0",x"20",x"11", -- 0x1168
		x"CD",x"E2",x"11",x"5F",x"78",x"07",x"CD",x"02", -- 0x1170
		x"11",x"3C",x"5A",x"CD",x"02",x"11",x"0D",x"18", -- 0x1178
		x"E5",x"67",x"E6",x"80",x"28",x"0F",x"5A",x"78", -- 0x1180
		x"C6",x"08",x"CD",x"02",x"11",x"7B",x"E6",x"10", -- 0x1188
		x"3E",x"0D",x"C4",x"02",x"11",x"7C",x"E6",x"40", -- 0x1190
		x"28",x"CC",x"CD",x"E2",x"11",x"57",x"CD",x"E2", -- 0x1198
		x"11",x"5F",x"3E",x"0B",x"CD",x"02",x"11",x"3C", -- 0x11A0
		x"5A",x"CD",x"02",x"11",x"0D",x"0D",x"18",x"B6", -- 0x11A8
		x"78",x"C6",x"08",x"1E",x"00",x"CD",x"02",x"11", -- 0x11B0
		x"04",x"21",x"3F",x"FB",x"AF",x"37",x"17",x"10", -- 0x11B8
		x"FD",x"A6",x"AE",x"77",x"3A",x"3F",x"FB",x"B7", -- 0x11C0
		x"C0",x"21",x"40",x"FB",x"7E",x"B7",x"C8",x"35", -- 0x11C8
		x"21",x"01",x"00",x"22",x"41",x"FB",x"22",x"66", -- 0x11D0
		x"FB",x"22",x"8B",x"FB",x"3E",x"07",x"32",x"3F", -- 0x11D8
		x"FB",x"C9",x"3A",x"3E",x"FB",x"E5",x"D5",x"C5", -- 0x11E0
		x"CD",x"AD",x"14",x"C3",x"DB",x"08",x"3D",x"FA", -- 0x11E8
		x"00",x"12",x"CD",x"0C",x"12",x"21",x"33",x"12", -- 0x11F0
		x"E6",x"0F",x"5F",x"16",x"00",x"19",x"7E",x"C9", -- 0x11F8
		x"CD",x"26",x"12",x"0F",x"0F",x"0F",x"0F",x"21", -- 0x1200
		x"43",x"12",x"18",x"EC",x"47",x"3E",x"0F",x"F3", -- 0x1208
		x"CD",x"0E",x"11",x"10",x"06",x"E6",x"DF",x"F6", -- 0x1210
		x"4C",x"18",x"04",x"E6",x"AF",x"F6",x"03",x"D3", -- 0x1218
		x"A1",x"CD",x"0C",x"11",x"FB",x"C9",x"F3",x"DB", -- 0x1220
		x"AA",x"E6",x"F0",x"C6",x"08",x"D3",x"AA",x"DB", -- 0x1228
		x"A9",x"FB",x"C9",x"00",x"05",x"01",x"00",x"03", -- 0x1230
		x"04",x"02",x"03",x"07",x"06",x"08",x"07",x"00", -- 0x1238
		x"05",x"01",x"00",x"00",x"03",x"05",x"04",x"01", -- 0x1240
		x"02",x"00",x"03",x"07",x"00",x"06",x"05",x"08", -- 0x1248
		x"01",x"07",x"00",x"3D",x"FA",x"6C",x"12",x"F5", -- 0x1250
		x"E6",x"01",x"CD",x"0C",x"12",x"C1",x"05",x"05", -- 0x1258
		x"06",x"10",x"FA",x"67",x"12",x"06",x"20",x"A0", -- 0x1260
		x"D6",x"01",x"9F",x"C9",x"CD",x"26",x"12",x"E6", -- 0x1268
		x"01",x"18",x"F5",x"3C",x"A7",x"1F",x"F5",x"47", -- 0x1270
		x"AF",x"37",x"17",x"10",x"FD",x"47",x"F1",x"0E", -- 0x1278
		x"10",x"11",x"AF",x"03",x"30",x"05",x"0E",x"20", -- 0x1280
		x"11",x"9F",x"4C",x"3E",x"0F",x"F3",x"CD",x"0E", -- 0x1288
		x"11",x"A3",x"B2",x"B1",x"D3",x"A1",x"A9",x"D3", -- 0x1290
		x"A1",x"3E",x"0E",x"D3",x"A0",x"0E",x"00",x"DB", -- 0x1298
		x"A2",x"A0",x"28",x"05",x"0C",x"C2",x"9F",x"12", -- 0x12A0
		x"0D",x"FB",x"79",x"C9",x"FE",x"04",x"11",x"EC", -- 0x12A8
		x"0C",x"38",x"05",x"11",x"D3",x"03",x"D6",x"04", -- 0x12B0
		x"3D",x"FA",x"C5",x"12",x"3D",x"3A",x"9D",x"FC", -- 0x12B8
		x"F8",x"3A",x"9C",x"FC",x"C8",x"F5",x"EB",x"22", -- 0x12C0
		x"66",x"F8",x"9F",x"2F",x"E6",x"40",x"4F",x"3E", -- 0x12C8
		x"0F",x"F3",x"CD",x"0E",x"11",x"E6",x"BF",x"B1", -- 0x12D0
		x"D3",x"A1",x"F1",x"FA",x"E8",x"12",x"CD",x"0C", -- 0x12D8
		x"11",x"FB",x"E6",x"08",x"D6",x"01",x"9F",x"C9", -- 0x12E0
		x"0E",x"00",x"CD",x"32",x"13",x"CD",x"32",x"13", -- 0x12E8
		x"38",x"28",x"CD",x"20",x"13",x"38",x"23",x"D5", -- 0x12F0
		x"CD",x"20",x"13",x"C1",x"38",x"1C",x"78",x"92", -- 0x12F8
		x"30",x"02",x"2F",x"3C",x"FE",x"05",x"30",x"E0", -- 0x1300
		x"79",x"93",x"30",x"02",x"2F",x"3C",x"FE",x"05", -- 0x1308
		x"30",x"D6",x"7A",x"32",x"9D",x"FC",x"7B",x"32", -- 0x1310
		x"9C",x"FC",x"FB",x"7C",x"D6",x"01",x"9F",x"C9", -- 0x1318
		x"0E",x"0A",x"CD",x"32",x"13",x"D8",x"55",x"D5", -- 0x1320
		x"0E",x"00",x"CD",x"32",x"13",x"D1",x"5D",x"AF", -- 0x1328
		x"67",x"C9",x"CD",x"5B",x"13",x"06",x"08",x"51", -- 0x1330
		x"CB",x"82",x"CB",x"92",x"CD",x"6D",x"13",x"CD", -- 0x1338
		x"0C",x"11",x"67",x"1F",x"1F",x"1F",x"CB",x"15", -- 0x1340
		x"CB",x"C2",x"CB",x"D2",x"CD",x"6D",x"13",x"10", -- 0x1348
		x"E7",x"CB",x"E2",x"CB",x"EA",x"CD",x"6D",x"13", -- 0x1350
		x"7C",x"1F",x"C9",x"3E",x"35",x"B1",x"57",x"CD", -- 0x1358
		x"6D",x"13",x"CD",x"0C",x"11",x"E6",x"02",x"28", -- 0x1360
		x"F9",x"CB",x"A2",x"CB",x"AA",x"E5",x"D5",x"2A", -- 0x1368
		x"66",x"F8",x"7D",x"2F",x"A2",x"57",x"3E",x"0F", -- 0x1370
		x"D3",x"A0",x"DB",x"A2",x"A5",x"B2",x"B4",x"D3", -- 0x1378
		x"A1",x"D1",x"E1",x"C9",x"A7",x"FA",x"92",x"13", -- 0x1380
		x"20",x"03",x"3E",x"09",x"C2",x"3E",x"08",x"D3", -- 0x1388
		x"AB",x"C9",x"DB",x"AA",x"E6",x"10",x"18",x"F0", -- 0x1390
		x"CD",x"D6",x"FD",x"ED",x"45",x"01",x"A0",x"00", -- 0x1398
		x"11",x"7F",x"F8",x"21",x"A9",x"13",x"ED",x"B0", -- 0x13A0
		x"C9",x"63",x"6F",x"6C",x"6F",x"72",x"20",x"00", -- 0x13A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13B0
		x"00",x"61",x"75",x"74",x"6F",x"20",x"00",x"00", -- 0x13B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13C0
		x"00",x"67",x"6F",x"74",x"6F",x"20",x"00",x"00", -- 0x13C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13D0
		x"00",x"6C",x"69",x"73",x"74",x"20",x"00",x"00", -- 0x13D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13E0
		x"00",x"72",x"75",x"6E",x"0D",x"00",x"00",x"00", -- 0x13E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13F0
		x"00",x"63",x"6F",x"6C",x"6F",x"72",x"20",x"31", -- 0x13F8
		x"35",x"2C",x"34",x"2C",x"34",x"0D",x"00",x"00", -- 0x1400
		x"00",x"63",x"6C",x"6F",x"61",x"64",x"22",x"00", -- 0x1408
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1410
		x"00",x"63",x"6F",x"6E",x"74",x"0D",x"00",x"00", -- 0x1418
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1420
		x"00",x"6C",x"69",x"73",x"74",x"2E",x"0D",x"1E", -- 0x1428
		x"1E",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1430
		x"00",x"0C",x"72",x"75",x"6E",x"0D",x"00",x"00", -- 0x1438
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1440
		x"00",x"DB",x"99",x"C9",x"DB",x"A8",x"C9",x"D3", -- 0x1448
		x"A8",x"C9",x"4F",x"F3",x"DB",x"AA",x"E6",x"F0", -- 0x1450
		x"81",x"D3",x"AA",x"DB",x"A9",x"FB",x"C9",x"CD", -- 0x1458
		x"DF",x"FE",x"E5",x"2A",x"64",x"F8",x"7D",x"B4", -- 0x1460
		x"E1",x"C9",x"7C",x"92",x"C0",x"7D",x"93",x"C9", -- 0x1468
		x"2E",x"02",x"18",x"03",x"3A",x"38",x"FB",x"D5", -- 0x1470
		x"11",x"41",x"FB",x"26",x"00",x"19",x"B7",x"28", -- 0x1478
		x"07",x"11",x"25",x"00",x"19",x"3D",x"20",x"FC", -- 0x1480
		x"D1",x"C9",x"CD",x"A7",x"FF",x"C9",x"CD",x"AC", -- 0x1488
		x"FF",x"C9",x"CD",x"FA",x"14",x"78",x"3C",x"23", -- 0x1490
		x"A6",x"B9",x"C8",x"E5",x"2B",x"2B",x"2B",x"E3", -- 0x1498
		x"23",x"4F",x"7E",x"23",x"66",x"6F",x"06",x"00", -- 0x14A0
		x"09",x"73",x"E1",x"71",x"C9",x"CD",x"FA",x"14", -- 0x14A8
		x"36",x"00",x"20",x"1D",x"79",x"B8",x"C8",x"23", -- 0x14B0
		x"3C",x"A6",x"2B",x"2B",x"E5",x"23",x"23",x"23", -- 0x14B8
		x"4F",x"7E",x"23",x"66",x"6F",x"06",x"00",x"09", -- 0x14C0
		x"7E",x"E1",x"71",x"B7",x"C0",x"3C",x"3E",x"00", -- 0x14C8
		x"C9",x"4F",x"06",x"00",x"21",x"70",x"F9",x"09", -- 0x14D0
		x"7E",x"C9",x"C5",x"CD",x"04",x"15",x"70",x"23", -- 0x14D8
		x"70",x"23",x"70",x"23",x"F1",x"77",x"23",x"73", -- 0x14E0
		x"23",x"72",x"C9",x"CD",x"FA",x"14",x"78",x"3C", -- 0x14E8
		x"23",x"A6",x"47",x"79",x"90",x"A6",x"6F",x"26", -- 0x14F0
		x"00",x"C9",x"CD",x"04",x"15",x"46",x"23",x"4E", -- 0x14F8
		x"23",x"7E",x"B7",x"C9",x"07",x"47",x"07",x"80", -- 0x1500
		x"4F",x"06",x"00",x"2A",x"F3",x"F3",x"09",x"C9", -- 0x1508
		x"E5",x"D5",x"C5",x"F5",x"CD",x"9D",x"08",x"30", -- 0x1510
		x"62",x"20",x"08",x"FE",x"0D",x"28",x"5F",x"FE", -- 0x1518
		x"20",x"38",x"58",x"CD",x"52",x"07",x"3A",x"E9", -- 0x1520
		x"F3",x"32",x"F2",x"F3",x"2A",x"B9",x"FC",x"EB", -- 0x1528
		x"ED",x"4B",x"B7",x"FC",x"CD",x"99",x"15",x"30", -- 0x1530
		x"42",x"CD",x"DF",x"15",x"11",x"40",x"FC",x"0E", -- 0x1538
		x"08",x"06",x"08",x"CD",x"39",x"16",x"E5",x"F5", -- 0x1540
		x"1A",x"87",x"F5",x"DC",x"7E",x"16",x"CD",x"AC", -- 0x1548
		x"16",x"E1",x"38",x"04",x"E5",x"F1",x"10",x"F1", -- 0x1550
		x"F1",x"E1",x"CD",x"40",x"16",x"CD",x"0A",x"17", -- 0x1558
		x"38",x"04",x"13",x"0D",x"20",x"DB",x"CD",x"D9", -- 0x1560
		x"15",x"3A",x"B7",x"FC",x"28",x"06",x"C6",x"20", -- 0x1568
		x"38",x"0C",x"18",x"04",x"C6",x"08",x"38",x"06", -- 0x1570
		x"32",x"B7",x"FC",x"C3",x"DA",x"08",x"AF",x"32", -- 0x1578
		x"B7",x"FC",x"CD",x"D9",x"15",x"3A",x"B9",x"FC", -- 0x1580
		x"28",x"03",x"C6",x"20",x"01",x"C6",x"08",x"FE", -- 0x1588
		x"C0",x"38",x"01",x"AF",x"32",x"B9",x"FC",x"18", -- 0x1590
		x"E2",x"E5",x"C5",x"06",x"01",x"EB",x"7C",x"87", -- 0x1598
		x"30",x"05",x"21",x"00",x"00",x"18",x"08",x"11", -- 0x15A0
		x"C0",x"00",x"E7",x"38",x"04",x"EB",x"2B",x"06", -- 0x15A8
		x"00",x"E3",x"7C",x"87",x"30",x"05",x"21",x"00", -- 0x15B0
		x"00",x"18",x"08",x"11",x"00",x"01",x"E7",x"38", -- 0x15B8
		x"04",x"EB",x"2B",x"06",x"00",x"D1",x"CD",x"D9", -- 0x15C0
		x"15",x"28",x"08",x"CB",x"3D",x"CB",x"3D",x"CB", -- 0x15C8
		x"3B",x"CB",x"3B",x"78",x"0F",x"44",x"4D",x"E1", -- 0x15D0
		x"C9",x"3A",x"AF",x"FC",x"D6",x"02",x"C9",x"C5", -- 0x15D8
		x"CD",x"D9",x"15",x"20",x"2E",x"51",x"79",x"E6", -- 0x15E0
		x"07",x"4F",x"21",x"0B",x"16",x"09",x"7E",x"32", -- 0x15E8
		x"2C",x"F9",x"7B",x"0F",x"0F",x"0F",x"E6",x"1F", -- 0x15F0
		x"47",x"7A",x"E6",x"F8",x"4F",x"7B",x"E6",x"07", -- 0x15F8
		x"B1",x"4F",x"2A",x"CB",x"F3",x"09",x"22",x"2A", -- 0x1600
		x"F9",x"C1",x"C9",x"80",x"40",x"20",x"10",x"08", -- 0x1608
		x"04",x"02",x"01",x"79",x"0F",x"3E",x"F0",x"30", -- 0x1610
		x"02",x"3E",x"0F",x"32",x"2C",x"F9",x"79",x"87", -- 0x1618
		x"87",x"E6",x"F8",x"4F",x"7B",x"E6",x"07",x"B1", -- 0x1620
		x"4F",x"7B",x"0F",x"0F",x"0F",x"E6",x"07",x"47", -- 0x1628
		x"2A",x"D5",x"F3",x"09",x"22",x"2A",x"F9",x"C1", -- 0x1630
		x"C9",x"3A",x"2C",x"F9",x"2A",x"2A",x"F9",x"C9", -- 0x1638
		x"32",x"2C",x"F9",x"22",x"2A",x"F9",x"C9",x"C5", -- 0x1640
		x"E5",x"CD",x"39",x"16",x"47",x"CD",x"D9",x"15", -- 0x1648
		x"20",x"1A",x"CD",x"D7",x"07",x"A0",x"F5",x"01", -- 0x1650
		x"00",x"20",x"09",x"CD",x"D7",x"07",x"47",x"F1", -- 0x1658
		x"78",x"28",x"04",x"0F",x"0F",x"0F",x"0F",x"E6", -- 0x1660
		x"0F",x"E1",x"C1",x"C9",x"CD",x"D7",x"07",x"04", -- 0x1668
		x"05",x"F2",x"67",x"16",x"18",x"ED",x"FE",x"10", -- 0x1670
		x"3F",x"D8",x"32",x"F2",x"F3",x"C9",x"E5",x"C5", -- 0x1678
		x"CD",x"D9",x"15",x"CD",x"39",x"16",x"20",x"08", -- 0x1680
		x"D5",x"CD",x"6C",x"18",x"D1",x"C1",x"E1",x"C9", -- 0x1688
		x"47",x"CD",x"D7",x"07",x"4F",x"78",x"2F",x"A1", -- 0x1690
		x"4F",x"3A",x"F2",x"F3",x"04",x"05",x"F2",x"A5", -- 0x1698
		x"16",x"87",x"87",x"87",x"87",x"B1",x"CD",x"CD", -- 0x16A0
		x"07",x"C1",x"E1",x"C9",x"E5",x"CD",x"D9",x"15", -- 0x16A8
		x"C2",x"79",x"17",x"CD",x"39",x"16",x"0F",x"30", -- 0x16B0
		x"4B",x"7D",x"E6",x"F8",x"FE",x"F8",x"3E",x"80", -- 0x16B8
		x"20",x"10",x"C3",x"5A",x"17",x"E5",x"CD",x"D9", -- 0x16C0
		x"15",x"C2",x"8B",x"17",x"CD",x"39",x"16",x"0F", -- 0x16C8
		x"30",x"32",x"D5",x"11",x"08",x"00",x"18",x"27", -- 0x16D0
		x"E5",x"CD",x"D9",x"15",x"C2",x"9C",x"17",x"CD", -- 0x16D8
		x"39",x"16",x"07",x"30",x"1F",x"7D",x"E6",x"F8", -- 0x16E0
		x"3E",x"01",x"20",x"0F",x"18",x"6C",x"E5",x"CD", -- 0x16E8
		x"D9",x"15",x"C2",x"AC",x"17",x"CD",x"39",x"16", -- 0x16F0
		x"07",x"30",x"09",x"D5",x"11",x"F8",x"FF",x"19", -- 0x16F8
		x"22",x"2A",x"F9",x"D1",x"32",x"2C",x"F9",x"A7", -- 0x1700
		x"E1",x"C9",x"E5",x"D5",x"2A",x"2A",x"F9",x"CD", -- 0x1708
		x"D9",x"15",x"C2",x"C6",x"17",x"E5",x"2A",x"CB", -- 0x1710
		x"F3",x"11",x"00",x"17",x"19",x"EB",x"E1",x"E7", -- 0x1718
		x"38",x"13",x"7D",x"3C",x"E6",x"07",x"20",x"0D", -- 0x1720
		x"18",x"2F",x"E5",x"D5",x"2A",x"2A",x"F9",x"CD", -- 0x1728
		x"D9",x"15",x"C2",x"DC",x"17",x"23",x"7D",x"11", -- 0x1730
		x"F8",x"00",x"18",x"31",x"E5",x"D5",x"2A",x"2A", -- 0x1738
		x"F9",x"CD",x"D9",x"15",x"C2",x"E3",x"17",x"E5", -- 0x1740
		x"2A",x"CB",x"F3",x"11",x"00",x"01",x"19",x"EB", -- 0x1748
		x"E1",x"E7",x"30",x"14",x"7D",x"E6",x"07",x"20", -- 0x1750
		x"0F",x"D1",x"37",x"E1",x"C9",x"E5",x"D5",x"2A", -- 0x1758
		x"2A",x"F9",x"CD",x"D9",x"15",x"C2",x"F8",x"17", -- 0x1760
		x"7D",x"2B",x"11",x"08",x"FF",x"E6",x"07",x"20", -- 0x1768
		x"01",x"19",x"22",x"2A",x"F9",x"A7",x"D1",x"E1", -- 0x1770
		x"C9",x"CD",x"39",x"16",x"A7",x"3E",x"0F",x"FA", -- 0x1778
		x"C0",x"17",x"7D",x"E6",x"F8",x"FE",x"F8",x"20", -- 0x1780
		x"0B",x"18",x"CF",x"CD",x"39",x"16",x"A7",x"3E", -- 0x1788
		x"0F",x"FA",x"C0",x"17",x"D5",x"11",x"08",x"00", -- 0x1790
		x"3E",x"F0",x"18",x"1F",x"CD",x"39",x"16",x"A7", -- 0x1798
		x"3E",x"F0",x"F2",x"C0",x"17",x"7D",x"E6",x"F8", -- 0x17A0
		x"20",x"0B",x"18",x"AE",x"CD",x"39",x"16",x"A7", -- 0x17A8
		x"3E",x"F0",x"F2",x"C0",x"17",x"D5",x"11",x"F8", -- 0x17B0
		x"FF",x"3E",x"0F",x"19",x"22",x"2A",x"F9",x"D1", -- 0x17B8
		x"32",x"2C",x"F9",x"A7",x"E1",x"C9",x"E5",x"2A", -- 0x17C0
		x"D5",x"F3",x"11",x"00",x"05",x"19",x"E1",x"E7", -- 0x17C8
		x"38",x"0A",x"7D",x"3C",x"E6",x"07",x"20",x"04", -- 0x17D0
		x"37",x"D1",x"E1",x"C9",x"23",x"7D",x"11",x"F8", -- 0x17D8
		x"00",x"18",x"1A",x"E5",x"2A",x"D5",x"F3",x"11", -- 0x17E0
		x"00",x"01",x"19",x"E1",x"E7",x"30",x"09",x"7D", -- 0x17E8
		x"E6",x"07",x"20",x"04",x"37",x"D1",x"E1",x"C9", -- 0x17F0
		x"7D",x"2B",x"11",x"08",x"FF",x"E6",x"07",x"20", -- 0x17F8
		x"01",x"19",x"22",x"2A",x"F9",x"A7",x"D1",x"E1", -- 0x1800
		x"C9",x"CD",x"D9",x"15",x"C2",x"BB",x"18",x"E5", -- 0x1808
		x"CD",x"39",x"16",x"E3",x"87",x"38",x"18",x"F5", -- 0x1810
		x"01",x"FF",x"FF",x"0F",x"09",x"30",x"45",x"0F", -- 0x1818
		x"30",x"FA",x"F1",x"3D",x"E3",x"E5",x"CD",x"6C", -- 0x1820
		x"18",x"E1",x"11",x"08",x"00",x"19",x"E3",x"7D", -- 0x1828
		x"E6",x"07",x"4F",x"7C",x"0F",x"7D",x"1F",x"0F", -- 0x1830
		x"0F",x"E6",x"3F",x"E1",x"47",x"28",x"14",x"AF", -- 0x1838
		x"CD",x"CD",x"07",x"11",x"00",x"20",x"19",x"3A", -- 0x1840
		x"F2",x"F3",x"CD",x"CD",x"07",x"11",x"08",x"20", -- 0x1848
		x"19",x"10",x"EC",x"0D",x"F8",x"E5",x"21",x"5D", -- 0x1850
		x"18",x"09",x"7E",x"18",x"0E",x"80",x"C0",x"E0", -- 0x1858
		x"F0",x"F8",x"FC",x"FE",x"87",x"3D",x"2F",x"47", -- 0x1860
		x"F1",x"3D",x"A0",x"E1",x"47",x"CD",x"D7",x"07", -- 0x1868
		x"4F",x"11",x"00",x"20",x"19",x"CD",x"D7",x"07", -- 0x1870
		x"F5",x"E6",x"0F",x"5F",x"F1",x"93",x"57",x"3A", -- 0x1878
		x"F2",x"F3",x"BB",x"28",x"19",x"87",x"87",x"87", -- 0x1880
		x"87",x"BA",x"28",x"16",x"F5",x"78",x"B1",x"FE", -- 0x1888
		x"FF",x"28",x"17",x"E5",x"D5",x"CD",x"A2",x"18", -- 0x1890
		x"D1",x"E1",x"F1",x"B3",x"18",x"1A",x"78",x"2F", -- 0x1898
		x"A1",x"11",x"78",x"B1",x"11",x"00",x"20",x"19", -- 0x18A0
		x"18",x"0E",x"F1",x"78",x"2F",x"E5",x"D5",x"CD", -- 0x18A8
		x"A4",x"18",x"D1",x"E1",x"3A",x"F2",x"F3",x"B2", -- 0x18B0
		x"C3",x"CD",x"07",x"E5",x"CD",x"7E",x"16",x"CD", -- 0x18B8
		x"C5",x"16",x"E1",x"2D",x"20",x"F5",x"C9",x"2A", -- 0x18C0
		x"0B",x"F4",x"EB",x"2A",x"0D",x"F4",x"C9",x"F5", -- 0x18C8
		x"CD",x"D9",x"15",x"28",x"06",x"F1",x"FE",x"10", -- 0x18D0
		x"3F",x"18",x"05",x"F1",x"3A",x"F2",x"F3",x"A7", -- 0x18D8
		x"32",x"B2",x"FC",x"C9",x"21",x"00",x"00",x"4D", -- 0x18E0
		x"CD",x"D9",x"15",x"20",x"64",x"78",x"32",x"66", -- 0x18E8
		x"F8",x"AF",x"32",x"69",x"F8",x"3A",x"B2",x"FC", -- 0x18F0
		x"47",x"CD",x"47",x"16",x"B8",x"20",x"0D",x"1B", -- 0x18F8
		x"7A",x"B3",x"C8",x"CD",x"AC",x"16",x"30",x"F1", -- 0x1900
		x"11",x"00",x"00",x"C9",x"CD",x"AE",x"19",x"D5", -- 0x1908
		x"CD",x"39",x"16",x"22",x"42",x"F9",x"32",x"44", -- 0x1910
		x"F9",x"11",x"00",x"00",x"13",x"CD",x"AC",x"16", -- 0x1918
		x"38",x"0B",x"CD",x"47",x"16",x"B8",x"28",x"05", -- 0x1920
		x"CD",x"AE",x"19",x"18",x"EF",x"D5",x"CD",x"39", -- 0x1928
		x"16",x"E5",x"F5",x"2A",x"42",x"F9",x"3A",x"44", -- 0x1930
		x"F9",x"CD",x"40",x"16",x"EB",x"22",x"67",x"F8", -- 0x1938
		x"3A",x"66",x"F8",x"A7",x"C4",x"09",x"18",x"F1", -- 0x1940
		x"E1",x"CD",x"40",x"16",x"E1",x"D1",x"C3",x"A9", -- 0x1948
		x"19",x"CD",x"C7",x"19",x"30",x"0D",x"1B",x"7A", -- 0x1950
		x"B3",x"C8",x"CD",x"AC",x"16",x"30",x"F2",x"11", -- 0x1958
		x"00",x"00",x"C9",x"CD",x"39",x"16",x"22",x"42", -- 0x1960
		x"F9",x"32",x"44",x"F9",x"21",x"00",x"00",x"23", -- 0x1968
		x"CD",x"AC",x"16",x"D8",x"CD",x"C7",x"19",x"30", -- 0x1970
		x"F6",x"C9",x"21",x"00",x"00",x"4D",x"CD",x"D9", -- 0x1978
		x"15",x"20",x"37",x"AF",x"32",x"69",x"F8",x"3A", -- 0x1980
		x"B2",x"FC",x"47",x"CD",x"D8",x"16",x"38",x"0F", -- 0x1988
		x"CD",x"47",x"16",x"B8",x"28",x"06",x"CD",x"AE", -- 0x1990
		x"19",x"23",x"18",x"EF",x"CD",x"C5",x"16",x"E5", -- 0x1998
		x"ED",x"5B",x"67",x"F8",x"19",x"CD",x"09",x"18", -- 0x19A0
		x"E1",x"3A",x"69",x"F8",x"4F",x"C9",x"E5",x"21", -- 0x19A8
		x"F2",x"F3",x"BE",x"E1",x"C8",x"3C",x"32",x"69", -- 0x19B0
		x"F8",x"C9",x"CD",x"D8",x"16",x"D8",x"CD",x"C7", -- 0x19B8
		x"19",x"DA",x"C5",x"16",x"23",x"18",x"F3",x"CD", -- 0x19C0
		x"47",x"16",x"47",x"3A",x"B2",x"FC",x"90",x"37", -- 0x19C8
		x"C8",x"3A",x"F2",x"F3",x"B8",x"C8",x"CD",x"7E", -- 0x19D0
		x"16",x"0E",x"01",x"A7",x"C9",x"C5",x"F5",x"01", -- 0x19D8
		x"00",x"00",x"0B",x"78",x"B1",x"20",x"FB",x"F1", -- 0x19E0
		x"C1",x"F5",x"3E",x"09",x"D3",x"AB",x"F1",x"FB", -- 0x19E8
		x"C9",x"B7",x"F5",x"3E",x"08",x"D3",x"AB",x"21", -- 0x19F0
		x"00",x"00",x"2B",x"7C",x"B5",x"20",x"FB",x"F1", -- 0x19F8
		x"3A",x"0A",x"F4",x"28",x"02",x"87",x"87",x"47", -- 0x1A00
		x"0E",x"00",x"F3",x"CD",x"4D",x"1A",x"CD",x"3F", -- 0x1A08
		x"1A",x"0B",x"78",x"B1",x"20",x"F5",x"C3",x"6F", -- 0x1A10
		x"04",x"2A",x"06",x"F4",x"F5",x"7D",x"D6",x"0E", -- 0x1A18
		x"6F",x"CD",x"50",x"1A",x"F1",x"06",x"08",x"0F", -- 0x1A20
		x"DC",x"40",x"1A",x"D4",x"39",x"1A",x"10",x"F7", -- 0x1A28
		x"CD",x"40",x"1A",x"CD",x"40",x"1A",x"C3",x"6F", -- 0x1A30
		x"04",x"2A",x"06",x"F4",x"CD",x"50",x"1A",x"C9", -- 0x1A38
		x"CD",x"4D",x"1A",x"E3",x"E3",x"00",x"00",x"00", -- 0x1A40
		x"00",x"CD",x"4D",x"1A",x"C9",x"2A",x"08",x"F4", -- 0x1A48
		x"F5",x"2D",x"C2",x"51",x"1A",x"3E",x"0B",x"D3", -- 0x1A50
		x"AB",x"25",x"C2",x"59",x"1A",x"3E",x"0A",x"D3", -- 0x1A58
		x"AB",x"F1",x"C9",x"3E",x"08",x"D3",x"AB",x"F3", -- 0x1A60
		x"3E",x"0E",x"D3",x"A0",x"21",x"57",x"04",x"51", -- 0x1A68
		x"CD",x"34",x"1B",x"D8",x"79",x"FE",x"DE",x"30", -- 0x1A70
		x"F3",x"FE",x"05",x"38",x"EF",x"92",x"30",x"02", -- 0x1A78
		x"2F",x"3C",x"FE",x"04",x"30",x"E6",x"2B",x"7C", -- 0x1A80
		x"B5",x"20",x"E4",x"21",x"00",x"00",x"45",x"55", -- 0x1A88
		x"CD",x"34",x"1B",x"D8",x"09",x"15",x"C2",x"90", -- 0x1A90
		x"1A",x"01",x"AE",x"06",x"09",x"7C",x"1F",x"E6", -- 0x1A98
		x"7F",x"57",x"29",x"7C",x"92",x"57",x"D6",x"06", -- 0x1AA0
		x"32",x"A4",x"FC",x"7A",x"87",x"06",x"00",x"D6", -- 0x1AA8
		x"03",x"04",x"30",x"FB",x"78",x"D6",x"03",x"32", -- 0x1AB0
		x"A5",x"FC",x"B7",x"C9",x"3A",x"A4",x"FC",x"57", -- 0x1AB8
		x"CD",x"6F",x"04",x"D8",x"DB",x"A2",x"07",x"30", -- 0x1AC0
		x"F7",x"CD",x"6F",x"04",x"D8",x"DB",x"A2",x"07", -- 0x1AC8
		x"38",x"F7",x"1E",x"00",x"CD",x"1F",x"1B",x"41", -- 0x1AD0
		x"CD",x"1F",x"1B",x"D8",x"78",x"81",x"DA",x"D7", -- 0x1AD8
		x"1A",x"BA",x"38",x"F3",x"2E",x"08",x"CD",x"03", -- 0x1AE0
		x"1B",x"FE",x"04",x"3F",x"D8",x"FE",x"02",x"3F", -- 0x1AE8
		x"CB",x"1A",x"79",x"0F",x"D4",x"23",x"1B",x"CD", -- 0x1AF0
		x"1F",x"1B",x"2D",x"C2",x"E6",x"1A",x"CD",x"6F", -- 0x1AF8
		x"04",x"7A",x"C9",x"3A",x"A5",x"FC",x"47",x"0E", -- 0x1B00
		x"00",x"DB",x"A2",x"AB",x"F2",x"17",x"1B",x"7B", -- 0x1B08
		x"2F",x"5F",x"0C",x"10",x"F4",x"79",x"C9",x"00", -- 0x1B10
		x"00",x"00",x"00",x"10",x"EC",x"79",x"C9",x"CD", -- 0x1B18
		x"6F",x"04",x"D8",x"0E",x"00",x"0C",x"28",x"0A", -- 0x1B20
		x"DB",x"A2",x"AB",x"F2",x"25",x"1B",x"7B",x"2F", -- 0x1B28
		x"5F",x"C9",x"0D",x"C9",x"CD",x"6F",x"04",x"D8", -- 0x1B30
		x"DB",x"A2",x"07",x"38",x"F7",x"1E",x"00",x"CD", -- 0x1B38
		x"23",x"1B",x"C3",x"25",x"1B",x"F5",x"CD",x"E4", -- 0x1B40
		x"FE",x"CD",x"5F",x"14",x"28",x"08",x"F1",x"DD", -- 0x1B48
		x"21",x"48",x"6C",x"C3",x"FF",x"01",x"3A",x"16", -- 0x1B50
		x"F4",x"B7",x"28",x"5F",x"3A",x"18",x"F4",x"A7", -- 0x1B58
		x"20",x"49",x"F1",x"F5",x"FE",x"09",x"20",x"0E", -- 0x1B60
		x"3E",x"20",x"CD",x"63",x"1B",x"3A",x"15",x"F4", -- 0x1B68
		x"E6",x"07",x"20",x"F4",x"F1",x"C9",x"D6",x"0D", -- 0x1B70
		x"28",x"0A",x"38",x"0B",x"FE",x"13",x"38",x"07", -- 0x1B78
		x"3A",x"15",x"F4",x"3C",x"32",x"15",x"F4",x"3A", -- 0x1B80
		x"17",x"F4",x"A7",x"28",x"1E",x"F1",x"CD",x"9D", -- 0x1B88
		x"08",x"D0",x"20",x"23",x"18",x"16",x"30",x"83", -- 0x1B90
		x"33",x"10",x"34",x"36",x"35",x"10",x"3A",x"C3", -- 0x1B98
		x"3C",x"10",x"3D",x"46",x"41",x"10",x"42",x"06", -- 0x1BA0
		x"FF",x"10",x"00",x"F1",x"CD",x"5D",x"08",x"D0", -- 0x1BA8
		x"DD",x"21",x"B2",x"73",x"C3",x"FF",x"01",x"3E", -- 0x1BB0
		x"20",x"18",x"F1",x"F1",x"C3",x"BC",x"08",x"00", -- 0x1BB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3C", -- 0x1BC0
		x"42",x"A5",x"81",x"A5",x"99",x"42",x"3C",x"3C", -- 0x1BC8
		x"7E",x"DB",x"FF",x"FF",x"DB",x"66",x"3C",x"6C", -- 0x1BD0
		x"FE",x"FE",x"FE",x"7C",x"38",x"10",x"00",x"10", -- 0x1BD8
		x"38",x"7C",x"FE",x"7C",x"38",x"10",x"00",x"10", -- 0x1BE0
		x"38",x"54",x"FE",x"54",x"10",x"38",x"00",x"10", -- 0x1BE8
		x"38",x"7C",x"FE",x"FE",x"10",x"38",x"00",x"00", -- 0x1BF0
		x"00",x"00",x"30",x"30",x"00",x"00",x"00",x"FF", -- 0x1BF8
		x"FF",x"FF",x"E7",x"E7",x"FF",x"FF",x"FF",x"38", -- 0x1C00
		x"44",x"82",x"82",x"82",x"44",x"38",x"00",x"C7", -- 0x1C08
		x"BB",x"7D",x"7D",x"7D",x"BB",x"C7",x"FF",x"0F", -- 0x1C10
		x"03",x"05",x"79",x"88",x"88",x"88",x"70",x"38", -- 0x1C18
		x"44",x"44",x"44",x"38",x"10",x"7C",x"10",x"30", -- 0x1C20
		x"28",x"24",x"24",x"28",x"20",x"E0",x"C0",x"3C", -- 0x1C28
		x"24",x"3C",x"24",x"24",x"E4",x"DC",x"18",x"10", -- 0x1C30
		x"54",x"38",x"EE",x"38",x"54",x"10",x"00",x"10", -- 0x1C38
		x"10",x"10",x"7C",x"10",x"10",x"10",x"10",x"10", -- 0x1C40
		x"10",x"10",x"FF",x"00",x"00",x"00",x"00",x"00", -- 0x1C48
		x"00",x"00",x"FF",x"10",x"10",x"10",x"10",x"10", -- 0x1C50
		x"10",x"10",x"F0",x"10",x"10",x"10",x"10",x"10", -- 0x1C58
		x"10",x"10",x"1F",x"10",x"10",x"10",x"10",x"10", -- 0x1C60
		x"10",x"10",x"FF",x"10",x"10",x"10",x"10",x"10", -- 0x1C68
		x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00", -- 0x1C70
		x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00", -- 0x1C78
		x"00",x"00",x"1F",x"10",x"10",x"10",x"10",x"00", -- 0x1C80
		x"00",x"00",x"F0",x"10",x"10",x"10",x"10",x"10", -- 0x1C88
		x"10",x"10",x"1F",x"00",x"00",x"00",x"00",x"10", -- 0x1C90
		x"10",x"10",x"F0",x"00",x"00",x"00",x"00",x"81", -- 0x1C98
		x"42",x"24",x"18",x"18",x"24",x"42",x"81",x"01", -- 0x1CA0
		x"02",x"04",x"08",x"10",x"20",x"40",x"80",x"80", -- 0x1CA8
		x"40",x"20",x"10",x"08",x"04",x"02",x"01",x"00", -- 0x1CB0
		x"10",x"10",x"FF",x"10",x"10",x"00",x"00",x"00", -- 0x1CB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20", -- 0x1CC0
		x"20",x"20",x"20",x"00",x"00",x"20",x"00",x"50", -- 0x1CC8
		x"50",x"50",x"00",x"00",x"00",x"00",x"00",x"50", -- 0x1CD0
		x"50",x"F8",x"50",x"F8",x"50",x"50",x"00",x"20", -- 0x1CD8
		x"78",x"A0",x"70",x"28",x"F0",x"20",x"00",x"C0", -- 0x1CE0
		x"C8",x"10",x"20",x"40",x"98",x"18",x"00",x"40", -- 0x1CE8
		x"A0",x"40",x"A8",x"90",x"98",x"60",x"00",x"10", -- 0x1CF0
		x"20",x"40",x"00",x"00",x"00",x"00",x"00",x"10", -- 0x1CF8
		x"20",x"40",x"40",x"40",x"20",x"10",x"00",x"40", -- 0x1D00
		x"20",x"10",x"10",x"10",x"20",x"40",x"00",x"20", -- 0x1D08
		x"A8",x"70",x"20",x"70",x"A8",x"20",x"00",x"00", -- 0x1D10
		x"20",x"20",x"F8",x"20",x"20",x"00",x"00",x"00", -- 0x1D18
		x"00",x"00",x"00",x"00",x"20",x"20",x"40",x"00", -- 0x1D20
		x"00",x"00",x"78",x"00",x"00",x"00",x"00",x"00", -- 0x1D28
		x"00",x"00",x"00",x"00",x"60",x"60",x"00",x"00", -- 0x1D30
		x"00",x"08",x"10",x"20",x"40",x"80",x"00",x"70", -- 0x1D38
		x"88",x"98",x"A8",x"C8",x"88",x"70",x"00",x"20", -- 0x1D40
		x"60",x"A0",x"20",x"20",x"20",x"F8",x"00",x"70", -- 0x1D48
		x"88",x"08",x"10",x"60",x"80",x"F8",x"00",x"70", -- 0x1D50
		x"88",x"08",x"30",x"08",x"88",x"70",x"00",x"10", -- 0x1D58
		x"30",x"50",x"90",x"F8",x"10",x"10",x"00",x"F8", -- 0x1D60
		x"80",x"E0",x"10",x"08",x"10",x"E0",x"00",x"30", -- 0x1D68
		x"40",x"80",x"F0",x"88",x"88",x"70",x"00",x"F8", -- 0x1D70
		x"88",x"10",x"20",x"20",x"20",x"20",x"00",x"70", -- 0x1D78
		x"88",x"88",x"70",x"88",x"88",x"70",x"00",x"70", -- 0x1D80
		x"88",x"88",x"78",x"08",x"10",x"60",x"00",x"00", -- 0x1D88
		x"00",x"20",x"00",x"00",x"20",x"00",x"00",x"00", -- 0x1D90
		x"00",x"20",x"00",x"00",x"20",x"20",x"40",x"18", -- 0x1D98
		x"30",x"60",x"C0",x"60",x"30",x"18",x"00",x"00", -- 0x1DA0
		x"00",x"F8",x"00",x"F8",x"00",x"00",x"00",x"C0", -- 0x1DA8
		x"60",x"30",x"18",x"30",x"60",x"C0",x"00",x"70", -- 0x1DB0
		x"88",x"08",x"10",x"20",x"00",x"20",x"00",x"70", -- 0x1DB8
		x"88",x"08",x"68",x"A8",x"A8",x"70",x"00",x"20", -- 0x1DC0
		x"50",x"88",x"88",x"F8",x"88",x"88",x"00",x"F0", -- 0x1DC8
		x"48",x"48",x"70",x"48",x"48",x"F0",x"00",x"30", -- 0x1DD0
		x"48",x"80",x"80",x"80",x"48",x"30",x"00",x"E0", -- 0x1DD8
		x"50",x"48",x"48",x"48",x"50",x"E0",x"00",x"F8", -- 0x1DE0
		x"80",x"80",x"F0",x"80",x"80",x"F8",x"00",x"F8", -- 0x1DE8
		x"80",x"80",x"F0",x"80",x"80",x"80",x"00",x"70", -- 0x1DF0
		x"88",x"80",x"B8",x"88",x"88",x"70",x"00",x"88", -- 0x1DF8
		x"88",x"88",x"F8",x"88",x"88",x"88",x"00",x"70", -- 0x1E00
		x"20",x"20",x"20",x"20",x"20",x"70",x"00",x"38", -- 0x1E08
		x"10",x"10",x"10",x"90",x"90",x"60",x"00",x"88", -- 0x1E10
		x"90",x"A0",x"C0",x"A0",x"90",x"88",x"00",x"80", -- 0x1E18
		x"80",x"80",x"80",x"80",x"80",x"F8",x"00",x"88", -- 0x1E20
		x"D8",x"A8",x"A8",x"88",x"88",x"88",x"00",x"88", -- 0x1E28
		x"C8",x"C8",x"A8",x"98",x"98",x"88",x"00",x"70", -- 0x1E30
		x"88",x"88",x"88",x"88",x"88",x"70",x"00",x"F0", -- 0x1E38
		x"88",x"88",x"F0",x"80",x"80",x"80",x"00",x"70", -- 0x1E40
		x"88",x"88",x"88",x"A8",x"90",x"68",x"00",x"F0", -- 0x1E48
		x"88",x"88",x"F0",x"A0",x"90",x"88",x"00",x"70", -- 0x1E50
		x"88",x"80",x"70",x"08",x"88",x"70",x"00",x"F8", -- 0x1E58
		x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"88", -- 0x1E60
		x"88",x"88",x"88",x"88",x"88",x"70",x"00",x"88", -- 0x1E68
		x"88",x"88",x"88",x"50",x"50",x"20",x"00",x"88", -- 0x1E70
		x"88",x"88",x"A8",x"A8",x"D8",x"88",x"00",x"88", -- 0x1E78
		x"88",x"50",x"20",x"50",x"88",x"88",x"00",x"88", -- 0x1E80
		x"88",x"88",x"70",x"20",x"20",x"20",x"00",x"F8", -- 0x1E88
		x"08",x"10",x"20",x"40",x"80",x"F8",x"00",x"70", -- 0x1E90
		x"40",x"40",x"40",x"40",x"40",x"70",x"00",x"00", -- 0x1E98
		x"00",x"80",x"40",x"20",x"10",x"08",x"00",x"70", -- 0x1EA0
		x"10",x"10",x"10",x"10",x"10",x"70",x"00",x"20", -- 0x1EA8
		x"50",x"88",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EB0
		x"00",x"00",x"00",x"00",x"00",x"F8",x"00",x"40", -- 0x1EB8
		x"20",x"10",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EC0
		x"00",x"70",x"08",x"78",x"88",x"78",x"00",x"80", -- 0x1EC8
		x"80",x"B0",x"C8",x"88",x"C8",x"B0",x"00",x"00", -- 0x1ED0
		x"00",x"70",x"88",x"80",x"88",x"70",x"00",x"08", -- 0x1ED8
		x"08",x"68",x"98",x"88",x"98",x"68",x"00",x"00", -- 0x1EE0
		x"00",x"70",x"88",x"F8",x"80",x"70",x"00",x"10", -- 0x1EE8
		x"28",x"20",x"F8",x"20",x"20",x"20",x"00",x"00", -- 0x1EF0
		x"00",x"68",x"98",x"98",x"68",x"08",x"70",x"80", -- 0x1EF8
		x"80",x"F0",x"88",x"88",x"88",x"88",x"00",x"20", -- 0x1F00
		x"00",x"60",x"20",x"20",x"20",x"70",x"00",x"10", -- 0x1F08
		x"00",x"30",x"10",x"10",x"10",x"90",x"60",x"40", -- 0x1F10
		x"40",x"48",x"50",x"60",x"50",x"48",x"00",x"60", -- 0x1F18
		x"20",x"20",x"20",x"20",x"20",x"70",x"00",x"00", -- 0x1F20
		x"00",x"D0",x"A8",x"A8",x"A8",x"A8",x"00",x"00", -- 0x1F28
		x"00",x"B0",x"C8",x"88",x"88",x"88",x"00",x"00", -- 0x1F30
		x"00",x"70",x"88",x"88",x"88",x"70",x"00",x"00", -- 0x1F38
		x"00",x"B0",x"C8",x"C8",x"B0",x"80",x"80",x"00", -- 0x1F40
		x"00",x"68",x"98",x"98",x"68",x"08",x"08",x"00", -- 0x1F48
		x"00",x"B0",x"C8",x"80",x"80",x"80",x"00",x"00", -- 0x1F50
		x"00",x"78",x"80",x"F0",x"08",x"F0",x"00",x"40", -- 0x1F58
		x"40",x"F0",x"40",x"40",x"48",x"30",x"00",x"00", -- 0x1F60
		x"00",x"90",x"90",x"90",x"90",x"68",x"00",x"00", -- 0x1F68
		x"00",x"88",x"88",x"88",x"50",x"20",x"00",x"00", -- 0x1F70
		x"00",x"88",x"A8",x"A8",x"A8",x"50",x"00",x"00", -- 0x1F78
		x"00",x"88",x"50",x"20",x"50",x"88",x"00",x"00", -- 0x1F80
		x"00",x"88",x"88",x"98",x"68",x"08",x"70",x"00", -- 0x1F88
		x"00",x"F8",x"10",x"20",x"40",x"F8",x"00",x"18", -- 0x1F90
		x"20",x"20",x"40",x"20",x"20",x"18",x"00",x"20", -- 0x1F98
		x"20",x"20",x"00",x"20",x"20",x"20",x"00",x"C0", -- 0x1FA0
		x"20",x"20",x"10",x"20",x"20",x"C0",x"00",x"40", -- 0x1FA8
		x"A8",x"10",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FB0
		x"00",x"20",x"50",x"F8",x"00",x"00",x"00",x"70", -- 0x1FB8
		x"88",x"80",x"80",x"88",x"70",x"20",x"60",x"90", -- 0x1FC0
		x"00",x"00",x"90",x"90",x"90",x"68",x"00",x"10", -- 0x1FC8
		x"20",x"70",x"88",x"F8",x"80",x"70",x"00",x"20", -- 0x1FD0
		x"50",x"70",x"08",x"78",x"88",x"78",x"00",x"48", -- 0x1FD8
		x"00",x"70",x"08",x"78",x"88",x"78",x"00",x"20", -- 0x1FE0
		x"10",x"70",x"08",x"78",x"88",x"78",x"00",x"20", -- 0x1FE8
		x"00",x"70",x"08",x"78",x"88",x"78",x"00",x"00", -- 0x1FF0
		x"70",x"80",x"80",x"80",x"70",x"10",x"60",x"20", -- 0x1FF8
		x"50",x"70",x"88",x"F8",x"80",x"70",x"00",x"50", -- 0x2000
		x"00",x"70",x"88",x"F8",x"80",x"70",x"00",x"20", -- 0x2008
		x"10",x"70",x"88",x"F8",x"80",x"70",x"00",x"50", -- 0x2010
		x"00",x"00",x"60",x"20",x"20",x"70",x"00",x"20", -- 0x2018
		x"50",x"00",x"60",x"20",x"20",x"70",x"00",x"40", -- 0x2020
		x"20",x"00",x"60",x"20",x"20",x"70",x"00",x"50", -- 0x2028
		x"00",x"20",x"50",x"88",x"F8",x"88",x"00",x"20", -- 0x2030
		x"00",x"20",x"50",x"88",x"F8",x"88",x"00",x"10", -- 0x2038
		x"20",x"F8",x"80",x"F0",x"80",x"F8",x"00",x"00", -- 0x2040
		x"00",x"6C",x"12",x"7E",x"90",x"6E",x"00",x"3E", -- 0x2048
		x"50",x"90",x"9C",x"F0",x"90",x"9E",x"00",x"60", -- 0x2050
		x"90",x"00",x"60",x"90",x"90",x"60",x"00",x"90", -- 0x2058
		x"00",x"00",x"60",x"90",x"90",x"60",x"00",x"40", -- 0x2060
		x"20",x"00",x"60",x"90",x"90",x"60",x"00",x"40", -- 0x2068
		x"A0",x"00",x"A0",x"A0",x"A0",x"50",x"00",x"40", -- 0x2070
		x"20",x"00",x"A0",x"A0",x"A0",x"50",x"00",x"90", -- 0x2078
		x"00",x"90",x"90",x"B0",x"50",x"10",x"E0",x"50", -- 0x2080
		x"00",x"70",x"88",x"88",x"88",x"70",x"00",x"50", -- 0x2088
		x"00",x"88",x"88",x"88",x"88",x"70",x"00",x"20", -- 0x2090
		x"20",x"78",x"80",x"80",x"78",x"20",x"20",x"18", -- 0x2098
		x"24",x"20",x"F8",x"20",x"E2",x"5C",x"00",x"88", -- 0x20A0
		x"50",x"20",x"F8",x"20",x"F8",x"20",x"00",x"C0", -- 0x20A8
		x"A0",x"A0",x"C8",x"9C",x"88",x"88",x"8C",x"18", -- 0x20B0
		x"20",x"20",x"F8",x"20",x"20",x"20",x"40",x"10", -- 0x20B8
		x"20",x"70",x"08",x"78",x"88",x"78",x"00",x"10", -- 0x20C0
		x"20",x"00",x"60",x"20",x"20",x"70",x"00",x"20", -- 0x20C8
		x"40",x"00",x"60",x"90",x"90",x"60",x"00",x"20", -- 0x20D0
		x"40",x"00",x"90",x"90",x"90",x"68",x"00",x"50", -- 0x20D8
		x"A0",x"00",x"A0",x"D0",x"90",x"90",x"00",x"28", -- 0x20E0
		x"50",x"00",x"C8",x"A8",x"98",x"88",x"00",x"00", -- 0x20E8
		x"70",x"08",x"78",x"88",x"78",x"00",x"F8",x"00", -- 0x20F0
		x"60",x"90",x"90",x"90",x"60",x"00",x"F0",x"20", -- 0x20F8
		x"00",x"20",x"40",x"80",x"88",x"70",x"00",x"00", -- 0x2100
		x"00",x"00",x"F8",x"80",x"80",x"00",x"00",x"00", -- 0x2108
		x"00",x"00",x"F8",x"08",x"08",x"00",x"00",x"84", -- 0x2110
		x"88",x"90",x"A8",x"54",x"84",x"08",x"1C",x"84", -- 0x2118
		x"88",x"90",x"A8",x"58",x"A8",x"3C",x"08",x"20", -- 0x2120
		x"00",x"00",x"20",x"20",x"20",x"20",x"00",x"00", -- 0x2128
		x"00",x"24",x"48",x"90",x"48",x"24",x"00",x"00", -- 0x2130
		x"00",x"90",x"48",x"24",x"48",x"90",x"00",x"28", -- 0x2138
		x"50",x"20",x"50",x"88",x"F8",x"88",x"00",x"28", -- 0x2140
		x"50",x"70",x"08",x"78",x"88",x"78",x"00",x"28", -- 0x2148
		x"50",x"00",x"70",x"20",x"20",x"70",x"00",x"28", -- 0x2150
		x"50",x"00",x"20",x"20",x"20",x"70",x"00",x"28", -- 0x2158
		x"50",x"00",x"70",x"88",x"88",x"70",x"00",x"50", -- 0x2160
		x"A0",x"00",x"60",x"90",x"90",x"60",x"00",x"28", -- 0x2168
		x"50",x"00",x"88",x"88",x"88",x"70",x"00",x"50", -- 0x2170
		x"A0",x"00",x"A0",x"A0",x"A0",x"50",x"00",x"FC", -- 0x2178
		x"48",x"48",x"48",x"E8",x"08",x"50",x"20",x"00", -- 0x2180
		x"50",x"00",x"50",x"50",x"50",x"10",x"20",x"C0", -- 0x2188
		x"44",x"C8",x"54",x"EC",x"54",x"9E",x"04",x"10", -- 0x2190
		x"A8",x"40",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2198
		x"20",x"50",x"88",x"50",x"20",x"00",x"00",x"88", -- 0x21A0
		x"10",x"20",x"40",x"80",x"28",x"00",x"00",x"7C", -- 0x21A8
		x"A8",x"A8",x"68",x"28",x"28",x"28",x"00",x"38", -- 0x21B0
		x"40",x"30",x"48",x"48",x"30",x"08",x"70",x"00", -- 0x21B8
		x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"F0", -- 0x21C0
		x"F0",x"F0",x"F0",x"0F",x"0F",x"0F",x"0F",x"00", -- 0x21C8
		x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x21D0
		x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x21D8
		x"00",x"00",x"3C",x"3C",x"00",x"00",x"00",x"FF", -- 0x21E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"C0", -- 0x21E8
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"0F", -- 0x21F0
		x"0F",x"0F",x"0F",x"F0",x"F0",x"F0",x"F0",x"FC", -- 0x21F8
		x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"03", -- 0x2200
		x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"3F", -- 0x2208
		x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"11", -- 0x2210
		x"22",x"44",x"88",x"11",x"22",x"44",x"88",x"88", -- 0x2218
		x"44",x"22",x"11",x"88",x"44",x"22",x"11",x"FE", -- 0x2220
		x"7C",x"38",x"10",x"00",x"00",x"00",x"00",x"00", -- 0x2228
		x"00",x"00",x"00",x"10",x"38",x"7C",x"FE",x"80", -- 0x2230
		x"C0",x"E0",x"F0",x"E0",x"C0",x"80",x"00",x"01", -- 0x2238
		x"03",x"07",x"0F",x"07",x"03",x"01",x"00",x"FF", -- 0x2240
		x"7E",x"3C",x"18",x"18",x"3C",x"7E",x"FF",x"81", -- 0x2248
		x"C3",x"E7",x"FF",x"FF",x"E7",x"C3",x"81",x"F0", -- 0x2250
		x"F0",x"F0",x"F0",x"00",x"00",x"00",x"00",x"00", -- 0x2258
		x"00",x"00",x"00",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x2260
		x"0F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"00", -- 0x2268
		x"00",x"00",x"00",x"F0",x"F0",x"F0",x"F0",x"33", -- 0x2270
		x"33",x"CC",x"CC",x"33",x"33",x"CC",x"CC",x"00", -- 0x2278
		x"20",x"20",x"50",x"50",x"88",x"F8",x"00",x"20", -- 0x2280
		x"20",x"70",x"20",x"70",x"20",x"20",x"00",x"00", -- 0x2288
		x"00",x"00",x"50",x"88",x"A8",x"50",x"00",x"FF", -- 0x2290
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00", -- 0x2298
		x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"F0", -- 0x22A0
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"0F", -- 0x22A8
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"FF", -- 0x22B0
		x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00", -- 0x22B8
		x"00",x"68",x"90",x"90",x"90",x"68",x"00",x"30", -- 0x22C0
		x"48",x"48",x"70",x"48",x"48",x"70",x"C0",x"F8", -- 0x22C8
		x"88",x"80",x"80",x"80",x"80",x"80",x"00",x"F8", -- 0x22D0
		x"50",x"50",x"50",x"50",x"50",x"98",x"00",x"F8", -- 0x22D8
		x"88",x"40",x"20",x"40",x"88",x"F8",x"00",x"00", -- 0x22E0
		x"00",x"78",x"90",x"90",x"90",x"60",x"00",x"00", -- 0x22E8
		x"50",x"50",x"50",x"50",x"68",x"80",x"80",x"00", -- 0x22F0
		x"50",x"A0",x"20",x"20",x"20",x"20",x"00",x"F8", -- 0x22F8
		x"20",x"70",x"A8",x"A8",x"70",x"20",x"F8",x"20", -- 0x2300
		x"50",x"88",x"F8",x"88",x"50",x"20",x"00",x"70", -- 0x2308
		x"88",x"88",x"88",x"50",x"50",x"D8",x"00",x"30", -- 0x2310
		x"40",x"40",x"20",x"50",x"50",x"50",x"20",x"00", -- 0x2318
		x"00",x"00",x"50",x"A8",x"A8",x"50",x"00",x"08", -- 0x2320
		x"70",x"A8",x"A8",x"A8",x"70",x"80",x"00",x"38", -- 0x2328
		x"40",x"80",x"F8",x"80",x"40",x"38",x"00",x"70", -- 0x2330
		x"88",x"88",x"88",x"88",x"88",x"88",x"00",x"00", -- 0x2338
		x"F8",x"00",x"F8",x"00",x"F8",x"00",x"00",x"20", -- 0x2340
		x"20",x"F8",x"20",x"20",x"00",x"F8",x"00",x"C0", -- 0x2348
		x"30",x"08",x"30",x"C0",x"00",x"F8",x"00",x"18", -- 0x2350
		x"60",x"80",x"60",x"18",x"00",x"F8",x"00",x"10", -- 0x2358
		x"28",x"20",x"20",x"20",x"20",x"20",x"20",x"20", -- 0x2360
		x"20",x"20",x"20",x"20",x"20",x"A0",x"40",x"00", -- 0x2368
		x"20",x"00",x"F8",x"00",x"20",x"00",x"00",x"00", -- 0x2370
		x"50",x"A0",x"00",x"50",x"A0",x"00",x"00",x"00", -- 0x2378
		x"18",x"24",x"24",x"18",x"00",x"00",x"00",x"00", -- 0x2380
		x"30",x"78",x"78",x"30",x"00",x"00",x"00",x"00", -- 0x2388
		x"00",x"00",x"00",x"30",x"00",x"00",x"00",x"3E", -- 0x2390
		x"20",x"20",x"20",x"A0",x"60",x"20",x"00",x"A0", -- 0x2398
		x"50",x"50",x"50",x"00",x"00",x"00",x"00",x"40", -- 0x23A0
		x"A0",x"20",x"40",x"E0",x"00",x"00",x"00",x"00", -- 0x23A8
		x"38",x"38",x"38",x"38",x"38",x"38",x"00",x"00", -- 0x23B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CD", -- 0x23B8
		x"DB",x"FD",x"3A",x"AA",x"F6",x"A7",x"20",x"0D", -- 0x23C0
		x"2E",x"00",x"18",x"14",x"CD",x"E0",x"FD",x"3E", -- 0x23C8
		x"3F",x"DF",x"3E",x"20",x"DF",x"CD",x"E5",x"FD", -- 0x23D0
		x"2A",x"DC",x"F3",x"2D",x"C4",x"29",x"0C",x"2C", -- 0x23D8
		x"22",x"CA",x"FB",x"AF",x"32",x"9B",x"FC",x"CD", -- 0x23E0
		x"CB",x"10",x"21",x"37",x"24",x"0E",x"0B",x"CD", -- 0x23E8
		x"19",x"09",x"F5",x"C4",x"FF",x"23",x"F1",x"30", -- 0x23F0
		x"EE",x"21",x"5D",x"F5",x"C8",x"3F",x"C9",x"F5", -- 0x23F8
		x"FE",x"09",x"20",x"0F",x"F1",x"3E",x"20",x"CD", -- 0x2400
		x"FF",x"23",x"3A",x"DD",x"F3",x"3D",x"E6",x"07", -- 0x2408
		x"20",x"F3",x"C9",x"F1",x"21",x"A8",x"FC",x"FE", -- 0x2410
		x"01",x"28",x"0B",x"FE",x"20",x"38",x"09",x"F5", -- 0x2418
		x"7E",x"A7",x"C4",x"F2",x"24",x"F1",x"DF",x"C9", -- 0x2420
		x"36",x"00",x"DF",x"3E",x"3E",x"AF",x"F5",x"CD", -- 0x2428
		x"2E",x"0A",x"F1",x"32",x"AA",x"FC",x"C3",x"E1", -- 0x2430
		x"09",x"08",x"61",x"25",x"12",x"E5",x"24",x"1B", -- 0x2438
		x"FE",x"23",x"02",x"0E",x"26",x"06",x"F8",x"25", -- 0x2440
		x"0E",x"D7",x"25",x"05",x"B9",x"25",x"03",x"C5", -- 0x2448
		x"24",x"0D",x"5A",x"24",x"15",x"AE",x"25",x"7F", -- 0x2450
		x"50",x"25",x"CD",x"6C",x"26",x"3A",x"AA",x"F6", -- 0x2458
		x"A7",x"28",x"02",x"26",x"01",x"E5",x"CD",x"2E", -- 0x2460
		x"0A",x"E1",x"11",x"5E",x"F5",x"06",x"FE",x"2D", -- 0x2468
		x"2C",x"D5",x"C5",x"CD",x"D8",x"0B",x"C1",x"D1", -- 0x2470
		x"A7",x"28",x"14",x"FE",x"20",x"30",x"0B",x"05", -- 0x2478
		x"28",x"1D",x"4F",x"3E",x"01",x"12",x"13",x"79", -- 0x2480
		x"C6",x"40",x"12",x"13",x"05",x"28",x"10",x"24", -- 0x2488
		x"3A",x"B0",x"F3",x"BC",x"30",x"DB",x"D5",x"CD", -- 0x2490
		x"1D",x"0C",x"D1",x"26",x"01",x"28",x"D1",x"1B", -- 0x2498
		x"1A",x"FE",x"20",x"28",x"FA",x"E5",x"D5",x"CD", -- 0x24A0
		x"E1",x"09",x"D1",x"E1",x"13",x"AF",x"12",x"3E", -- 0x24A8
		x"0D",x"A7",x"F5",x"CD",x"29",x"0C",x"CD",x"8E", -- 0x24B0
		x"08",x"3E",x"0A",x"DF",x"AF",x"32",x"A8",x"FC", -- 0x24B8
		x"F1",x"37",x"E1",x"C9",x"2C",x"CD",x"1D",x"0C", -- 0x24C0
		x"28",x"FA",x"CD",x"2D",x"24",x"AF",x"32",x"5E", -- 0x24C8
		x"F5",x"26",x"01",x"E5",x"CD",x"BD",x"04",x"CD", -- 0x24D0
		x"54",x"04",x"E1",x"38",x"D2",x"3A",x"B1",x"FB", -- 0x24D8
		x"A7",x"20",x"CC",x"18",x"CD",x"21",x"A8",x"FC", -- 0x24E0
		x"7E",x"EE",x"FF",x"77",x"CA",x"2D",x"24",x"C3", -- 0x24E8
		x"2C",x"24",x"CD",x"2E",x"0A",x"2A",x"DC",x"F3", -- 0x24F0
		x"0E",x"20",x"E5",x"C5",x"CD",x"D8",x"0B",x"D1", -- 0x24F8
		x"C5",x"4B",x"CD",x"E6",x"0B",x"C1",x"3A",x"B0", -- 0x2500
		x"F3",x"24",x"BC",x"7A",x"30",x"ED",x"E1",x"CD", -- 0x2508
		x"1D",x"0C",x"28",x"37",x"79",x"FE",x"20",x"F5", -- 0x2510
		x"20",x"0A",x"3A",x"B0",x"F3",x"BC",x"28",x"04", -- 0x2518
		x"F1",x"C3",x"E1",x"09",x"CD",x"2A",x"0C",x"2C", -- 0x2520
		x"C5",x"E5",x"CD",x"32",x"0C",x"BD",x"38",x"05", -- 0x2528
		x"CD",x"B7",x"0A",x"18",x"0F",x"21",x"DC",x"F3", -- 0x2530
		x"35",x"20",x"01",x"34",x"2E",x"01",x"CD",x"88", -- 0x2538
		x"0A",x"E1",x"2D",x"E5",x"E1",x"C1",x"F1",x"CA", -- 0x2540
		x"E1",x"09",x"2D",x"2C",x"26",x"01",x"18",x"AA", -- 0x2548
		x"3A",x"B0",x"F3",x"BC",x"20",x"05",x"CD",x"1D", -- 0x2550
		x"0C",x"20",x"3A",x"3E",x"1C",x"DF",x"2A",x"DC", -- 0x2558
		x"F3",x"E5",x"CD",x"2E",x"0A",x"E1",x"25",x"C2", -- 0x2560
		x"7A",x"25",x"24",x"E5",x"2D",x"28",x"0A",x"3A", -- 0x2568
		x"B0",x"F3",x"67",x"CD",x"1D",x"0C",x"20",x"01", -- 0x2570
		x"E3",x"E1",x"22",x"DC",x"F3",x"3A",x"B0",x"F3", -- 0x2578
		x"BC",x"28",x"12",x"24",x"CD",x"D8",x"0B",x"25", -- 0x2580
		x"CD",x"E6",x"0B",x"24",x"24",x"3A",x"B0",x"F3", -- 0x2588
		x"3C",x"BC",x"20",x"F0",x"25",x"0E",x"20",x"CD", -- 0x2590
		x"E6",x"0B",x"CD",x"1D",x"0C",x"C2",x"E1",x"09", -- 0x2598
		x"E5",x"2C",x"26",x"01",x"CD",x"D8",x"0B",x"E3", -- 0x25A0
		x"CD",x"E6",x"0B",x"E1",x"18",x"CF",x"CD",x"2E", -- 0x25A8
		x"0A",x"CD",x"6C",x"26",x"22",x"DC",x"F3",x"18", -- 0x25B0
		x"05",x"E5",x"CD",x"2E",x"0A",x"E1",x"CD",x"1D", -- 0x25B8
		x"0C",x"F5",x"CD",x"EE",x"0A",x"F1",x"20",x"05", -- 0x25C0
		x"26",x"01",x"2C",x"18",x"F1",x"CD",x"E1",x"09", -- 0x25C8
		x"AF",x"32",x"A8",x"FC",x"C3",x"2D",x"24",x"CD", -- 0x25D0
		x"2E",x"0A",x"2A",x"DC",x"F3",x"2D",x"2C",x"CD", -- 0x25D8
		x"1D",x"0C",x"28",x"FA",x"3A",x"B0",x"F3",x"67", -- 0x25E0
		x"24",x"25",x"28",x"07",x"CD",x"D8",x"0B",x"FE", -- 0x25E8
		x"20",x"28",x"F6",x"CD",x"5B",x"0A",x"18",x"D5", -- 0x25F0
		x"CD",x"2E",x"0A",x"CD",x"34",x"26",x"CD",x"24", -- 0x25F8
		x"26",x"28",x"CA",x"38",x"F9",x"CD",x"24",x"26", -- 0x2600
		x"28",x"C3",x"30",x"F9",x"18",x"BF",x"CD",x"2E", -- 0x2608
		x"0A",x"CD",x"34",x"26",x"28",x"B7",x"30",x"F9", -- 0x2610
		x"CD",x"34",x"26",x"28",x"B0",x"38",x"F9",x"CD", -- 0x2618
		x"5B",x"0A",x"18",x"A9",x"2A",x"DC",x"F3",x"CD", -- 0x2620
		x"5B",x"0A",x"CD",x"32",x"0C",x"5F",x"3A",x"B0", -- 0x2628
		x"F3",x"57",x"18",x"09",x"2A",x"DC",x"F3",x"CD", -- 0x2630
		x"4C",x"0A",x"11",x"01",x"01",x"2A",x"DC",x"F3", -- 0x2638
		x"E7",x"C8",x"11",x"68",x"26",x"D5",x"CD",x"D8", -- 0x2640
		x"0B",x"FE",x"30",x"3F",x"D0",x"FE",x"3A",x"D8", -- 0x2648
		x"FE",x"41",x"3F",x"D0",x"FE",x"5B",x"D8",x"FE", -- 0x2650
		x"61",x"3F",x"D0",x"FE",x"7B",x"D8",x"FE",x"86", -- 0x2658
		x"3F",x"D0",x"FE",x"A0",x"D8",x"FE",x"A6",x"3F", -- 0x2660
		x"3E",x"00",x"3C",x"C9",x"2D",x"28",x"05",x"CD", -- 0x2668
		x"1D",x"0C",x"28",x"F8",x"2C",x"3A",x"CA",x"FB", -- 0x2670
		x"BD",x"26",x"01",x"C0",x"2A",x"CA",x"FB",x"C9", -- 0x2678
		x"C3",x"76",x"7C",x"C3",x"8C",x"55",x"C3",x"66", -- 0x2680
		x"46",x"C3",x"97",x"55",x"21",x"47",x"F8",x"7E", -- 0x2688
		x"B7",x"C8",x"EE",x"80",x"77",x"18",x"09",x"CD", -- 0x2690
		x"EF",x"2E",x"21",x"47",x"F8",x"7E",x"B7",x"C8", -- 0x2698
		x"E6",x"7F",x"47",x"11",x"F6",x"F7",x"1A",x"B7", -- 0x26A0
		x"CA",x"05",x"2F",x"E6",x"7F",x"90",x"30",x"11", -- 0x26A8
		x"2F",x"3C",x"F5",x"E5",x"06",x"08",x"1A",x"4E", -- 0x26B0
		x"77",x"79",x"12",x"13",x"23",x"10",x"F7",x"E1", -- 0x26B8
		x"F1",x"FE",x"10",x"D0",x"F5",x"AF",x"32",x"FE", -- 0x26C0
		x"F7",x"32",x"4F",x"F8",x"21",x"48",x"F8",x"F1", -- 0x26C8
		x"CD",x"A3",x"27",x"21",x"47",x"F8",x"3A",x"F6", -- 0x26D0
		x"F7",x"AE",x"FA",x"F7",x"26",x"3A",x"4F",x"F8", -- 0x26D8
		x"32",x"FE",x"F7",x"CD",x"59",x"27",x"D2",x"3C", -- 0x26E0
		x"27",x"EB",x"7E",x"34",x"AE",x"FA",x"67",x"40", -- 0x26E8
		x"CD",x"DB",x"27",x"CB",x"E6",x"18",x"45",x"CD", -- 0x26F0
		x"6B",x"27",x"21",x"F7",x"F7",x"01",x"00",x"08", -- 0x26F8
		x"7E",x"B7",x"20",x"08",x"23",x"0D",x"0D",x"10", -- 0x2700
		x"F7",x"C3",x"7D",x"2E",x"E6",x"F0",x"20",x"06", -- 0x2708
		x"E5",x"CD",x"97",x"27",x"E1",x"0D",x"3E",x"08", -- 0x2710
		x"90",x"28",x"12",x"F5",x"C5",x"48",x"11",x"F7", -- 0x2718
		x"F7",x"06",x"00",x"ED",x"B0",x"C1",x"F1",x"47", -- 0x2720
		x"AF",x"12",x"13",x"10",x"FC",x"79",x"B7",x"28", -- 0x2728
		x"0B",x"21",x"F6",x"F7",x"46",x"86",x"77",x"A8", -- 0x2730
		x"FA",x"67",x"40",x"C8",x"21",x"FE",x"F7",x"06", -- 0x2738
		x"07",x"7E",x"FE",x"50",x"D8",x"2B",x"AF",x"37", -- 0x2740
		x"8E",x"27",x"77",x"D0",x"2B",x"10",x"F9",x"7E", -- 0x2748
		x"34",x"AE",x"FA",x"67",x"40",x"23",x"36",x"10", -- 0x2750
		x"C9",x"21",x"4E",x"F8",x"11",x"FD",x"F7",x"06", -- 0x2758
		x"07",x"AF",x"1A",x"8E",x"27",x"12",x"1B",x"2B", -- 0x2760
		x"10",x"F8",x"C9",x"21",x"4F",x"F8",x"7E",x"FE", -- 0x2768
		x"50",x"20",x"01",x"34",x"11",x"FE",x"F7",x"06", -- 0x2770
		x"08",x"AF",x"1A",x"9E",x"27",x"12",x"1B",x"2B", -- 0x2778
		x"10",x"F8",x"D0",x"EB",x"7E",x"EE",x"80",x"77", -- 0x2780
		x"21",x"FE",x"F7",x"06",x"08",x"AF",x"3E",x"00", -- 0x2788
		x"9E",x"27",x"77",x"2B",x"10",x"F8",x"C9",x"21", -- 0x2790
		x"FE",x"F7",x"C5",x"AF",x"ED",x"6F",x"2B",x"10", -- 0x2798
		x"FB",x"C1",x"C9",x"B7",x"1F",x"F5",x"B7",x"CA", -- 0x27A0
		x"E2",x"27",x"F5",x"2F",x"3C",x"4F",x"06",x"FF", -- 0x27A8
		x"11",x"07",x"00",x"19",x"54",x"5D",x"09",x"3E", -- 0x27B0
		x"08",x"81",x"4F",x"C5",x"06",x"00",x"ED",x"B8", -- 0x27B8
		x"C1",x"F1",x"23",x"13",x"D5",x"47",x"AF",x"77", -- 0x27C0
		x"23",x"10",x"FC",x"E1",x"F1",x"D0",x"79",x"E5", -- 0x27C8
		x"C5",x"47",x"AF",x"ED",x"67",x"23",x"10",x"FB", -- 0x27D0
		x"C1",x"E1",x"C9",x"21",x"F7",x"F7",x"3E",x"08", -- 0x27D8
		x"18",x"ED",x"F1",x"D0",x"18",x"F8",x"CD",x"71", -- 0x27E0
		x"2E",x"C8",x"3A",x"47",x"F8",x"B7",x"CA",x"7D", -- 0x27E8
		x"2E",x"47",x"21",x"F6",x"F7",x"AE",x"E6",x"80", -- 0x27F0
		x"4F",x"CB",x"B8",x"7E",x"E6",x"7F",x"80",x"47", -- 0x27F8
		x"36",x"00",x"E6",x"C0",x"C8",x"FE",x"C0",x"20", -- 0x2800
		x"03",x"C3",x"67",x"40",x"78",x"C6",x"40",x"E6", -- 0x2808
		x"7F",x"C8",x"B1",x"2B",x"77",x"11",x"45",x"F8", -- 0x2810
		x"01",x"08",x"00",x"21",x"FD",x"F7",x"D5",x"ED", -- 0x2818
		x"B8",x"23",x"AF",x"06",x"08",x"77",x"23",x"10", -- 0x2820
		x"FC",x"D1",x"01",x"83",x"28",x"C5",x"CD",x"8A", -- 0x2828
		x"28",x"E5",x"01",x"08",x"00",x"EB",x"ED",x"B8", -- 0x2830
		x"EB",x"21",x"3D",x"F8",x"06",x"08",x"CD",x"61", -- 0x2838
		x"27",x"D1",x"CD",x"8A",x"28",x"0E",x"07",x"11", -- 0x2840
		x"4E",x"F8",x"1A",x"B7",x"20",x"04",x"1B",x"0D", -- 0x2848
		x"18",x"F8",x"1A",x"1B",x"D5",x"21",x"0D",x"F8", -- 0x2850
		x"87",x"38",x"08",x"28",x"14",x"11",x"08",x"00", -- 0x2858
		x"19",x"18",x"F5",x"F5",x"06",x"08",x"11",x"FD", -- 0x2860
		x"F7",x"E5",x"CD",x"61",x"27",x"E1",x"F1",x"18", -- 0x2868
		x"EC",x"06",x"0F",x"11",x"04",x"F8",x"21",x"05", -- 0x2870
		x"F8",x"CD",x"FE",x"2E",x"36",x"00",x"D1",x"0D", -- 0x2878
		x"20",x"D0",x"C9",x"2B",x"7E",x"23",x"77",x"C3", -- 0x2880
		x"FA",x"26",x"21",x"F8",x"FF",x"19",x"0E",x"03", -- 0x2888
		x"06",x"08",x"B7",x"1A",x"8F",x"27",x"77",x"2B", -- 0x2890
		x"1B",x"10",x"F8",x"0D",x"20",x"F2",x"C9",x"3A", -- 0x2898
		x"47",x"F8",x"B7",x"CA",x"58",x"40",x"47",x"21", -- 0x28A0
		x"F6",x"F7",x"7E",x"B7",x"CA",x"7D",x"2E",x"A8", -- 0x28A8
		x"E6",x"80",x"4F",x"CB",x"B8",x"7E",x"E6",x"7F", -- 0x28B0
		x"90",x"47",x"1F",x"A8",x"E6",x"40",x"36",x"00", -- 0x28B8
		x"28",x"07",x"78",x"E6",x"80",x"C0",x"C3",x"67", -- 0x28C0
		x"40",x"78",x"C6",x"41",x"E6",x"7F",x"77",x"28", -- 0x28C8
		x"F5",x"B1",x"36",x"00",x"2B",x"77",x"11",x"FD", -- 0x28D0
		x"F7",x"21",x"4E",x"F8",x"06",x"07",x"AF",x"BE", -- 0x28D8
		x"20",x"04",x"1B",x"2B",x"10",x"F9",x"22",x"F2", -- 0x28E0
		x"F7",x"EB",x"22",x"F0",x"F7",x"78",x"32",x"F4", -- 0x28E8
		x"F7",x"21",x"3E",x"F8",x"06",x"0F",x"E5",x"C5", -- 0x28F0
		x"2A",x"F2",x"F7",x"EB",x"2A",x"F0",x"F7",x"3A", -- 0x28F8
		x"F4",x"F7",x"0E",x"FF",x"0C",x"47",x"E5",x"D5", -- 0x2900
		x"AF",x"EB",x"1A",x"9E",x"27",x"12",x"2B",x"1B", -- 0x2908
		x"10",x"F8",x"1A",x"98",x"12",x"D1",x"E1",x"3A", -- 0x2910
		x"F4",x"F7",x"30",x"E8",x"47",x"EB",x"CD",x"61", -- 0x2918
		x"27",x"30",x"02",x"EB",x"34",x"79",x"C1",x"4F", -- 0x2920
		x"C5",x"CB",x"38",x"04",x"58",x"16",x"00",x"21", -- 0x2928
		x"F5",x"F7",x"19",x"CD",x"9A",x"27",x"C1",x"E1", -- 0x2930
		x"78",x"0C",x"0D",x"20",x"36",x"FE",x"0F",x"28", -- 0x2938
		x"23",x"0F",x"07",x"30",x"2E",x"C5",x"E5",x"21", -- 0x2940
		x"F6",x"F7",x"06",x"08",x"AF",x"BE",x"20",x"0F", -- 0x2948
		x"23",x"10",x"FA",x"E1",x"C1",x"CB",x"38",x"04", -- 0x2950
		x"AF",x"77",x"23",x"10",x"FC",x"18",x"26",x"E1", -- 0x2958
		x"C1",x"78",x"18",x"0F",x"3A",x"F5",x"F7",x"5F", -- 0x2960
		x"3D",x"32",x"F5",x"F7",x"AB",x"F2",x"F4",x"28", -- 0x2968
		x"C3",x"7D",x"2E",x"1F",x"79",x"38",x"05",x"B6", -- 0x2970
		x"77",x"23",x"18",x"05",x"87",x"87",x"87",x"87", -- 0x2978
		x"77",x"05",x"C2",x"F6",x"28",x"21",x"FE",x"F7", -- 0x2980
		x"11",x"45",x"F8",x"06",x"08",x"CD",x"FE",x"2E", -- 0x2988
		x"C3",x"83",x"28",x"21",x"63",x"2D",x"CD",x"3B", -- 0x2990
		x"2C",x"3A",x"F6",x"F7",x"E6",x"7F",x"32",x"F6", -- 0x2998
		x"F7",x"21",x"23",x"2D",x"CD",x"32",x"2C",x"CD", -- 0x29A0
		x"8D",x"2E",x"18",x"06",x"21",x"63",x"2D",x"CD", -- 0x29A8
		x"3B",x"2C",x"3A",x"F6",x"F7",x"B7",x"FC",x"80", -- 0x29B0
		x"2C",x"CD",x"CC",x"2C",x"CD",x"CF",x"30",x"CD", -- 0x29B8
		x"4D",x"2C",x"CD",x"E1",x"2C",x"CD",x"8C",x"26", -- 0x29C0
		x"3A",x"F6",x"F7",x"FE",x"40",x"DA",x"F5",x"29", -- 0x29C8
		x"3A",x"F7",x"F7",x"FE",x"25",x"DA",x"F5",x"29", -- 0x29D0
		x"FE",x"75",x"D2",x"EC",x"29",x"CD",x"4D",x"2C", -- 0x29D8
		x"21",x"11",x"2D",x"CD",x"5C",x"2C",x"CD",x"8C", -- 0x29E0
		x"26",x"C3",x"F5",x"29",x"21",x"1B",x"2D",x"CD", -- 0x29E8
		x"50",x"2C",x"CD",x"8C",x"26",x"21",x"EF",x"2D", -- 0x29F0
		x"C3",x"88",x"2C",x"CD",x"CC",x"2C",x"CD",x"93", -- 0x29F8
		x"29",x"CD",x"6F",x"2C",x"CD",x"AC",x"29",x"CD", -- 0x2A00
		x"DC",x"2C",x"3A",x"47",x"F8",x"B7",x"C2",x"9F", -- 0x2A08
		x"28",x"C3",x"67",x"40",x"3A",x"F6",x"F7",x"B7", -- 0x2A10
		x"C8",x"FC",x"80",x"2C",x"FE",x"41",x"DA",x"3C", -- 0x2A18
		x"2A",x"CD",x"4D",x"2C",x"21",x"1B",x"2D",x"CD", -- 0x2A20
		x"5C",x"2C",x"CD",x"9F",x"28",x"CD",x"3C",x"2A", -- 0x2A28
		x"CD",x"4D",x"2C",x"21",x"43",x"2D",x"CD",x"5C", -- 0x2A30
		x"2C",x"C3",x"8C",x"26",x"21",x"4B",x"2D",x"CD", -- 0x2A38
		x"47",x"2C",x"FA",x"6C",x"2A",x"CD",x"CC",x"2C", -- 0x2A40
		x"21",x"53",x"2D",x"CD",x"2C",x"2C",x"CD",x"6F", -- 0x2A48
		x"2C",x"21",x"53",x"2D",x"CD",x"3B",x"2C",x"21", -- 0x2A50
		x"1B",x"2D",x"CD",x"32",x"2C",x"CD",x"DC",x"2C", -- 0x2A58
		x"CD",x"9F",x"28",x"CD",x"6C",x"2A",x"21",x"5B", -- 0x2A60
		x"2D",x"C3",x"2C",x"2C",x"21",x"30",x"2E",x"C3", -- 0x2A68
		x"88",x"2C",x"CD",x"71",x"2E",x"FA",x"5A",x"47", -- 0x2A70
		x"CA",x"5A",x"47",x"21",x"F6",x"F7",x"7E",x"F5", -- 0x2A78
		x"36",x"41",x"21",x"2B",x"2D",x"CD",x"47",x"2C", -- 0x2A80
		x"FA",x"92",x"2A",x"F1",x"3C",x"F5",x"21",x"F6", -- 0x2A88
		x"F7",x"35",x"F1",x"32",x"9D",x"F6",x"CD",x"CC", -- 0x2A90
		x"2C",x"21",x"1B",x"2D",x"CD",x"2C",x"2C",x"CD", -- 0x2A98
		x"6F",x"2C",x"21",x"1B",x"2D",x"CD",x"32",x"2C", -- 0x2AA0
		x"CD",x"DC",x"2C",x"CD",x"9F",x"28",x"CD",x"CC", -- 0x2AA8
		x"2C",x"CD",x"38",x"2C",x"CD",x"CC",x"2C",x"CD", -- 0x2AB0
		x"CC",x"2C",x"21",x"C6",x"2D",x"CD",x"A3",x"2C", -- 0x2AB8
		x"CD",x"6F",x"2C",x"21",x"A5",x"2D",x"CD",x"A3", -- 0x2AC0
		x"2C",x"CD",x"DC",x"2C",x"CD",x"9F",x"28",x"CD", -- 0x2AC8
		x"DC",x"2C",x"CD",x"E6",x"27",x"21",x"33",x"2D", -- 0x2AD0
		x"CD",x"2C",x"2C",x"CD",x"DC",x"2C",x"CD",x"E6", -- 0x2AD8
		x"27",x"CD",x"CC",x"2C",x"3A",x"9D",x"F6",x"D6", -- 0x2AE0
		x"41",x"6F",x"87",x"9F",x"67",x"CD",x"CB",x"2F", -- 0x2AE8
		x"CD",x"42",x"30",x"CD",x"DC",x"2C",x"CD",x"9A", -- 0x2AF0
		x"26",x"21",x"3B",x"2D",x"C3",x"3B",x"2C",x"CD", -- 0x2AF8
		x"71",x"2E",x"C8",x"FA",x"5A",x"47",x"CD",x"4D", -- 0x2B00
		x"2C",x"3A",x"F6",x"F7",x"B7",x"1F",x"CE",x"20", -- 0x2B08
		x"32",x"47",x"F8",x"3A",x"F7",x"F7",x"B7",x"0F", -- 0x2B10
		x"B7",x"0F",x"E6",x"33",x"C6",x"10",x"32",x"48", -- 0x2B18
		x"F8",x"3E",x"07",x"32",x"9D",x"F6",x"CD",x"CC", -- 0x2B20
		x"2C",x"CD",x"C7",x"2C",x"CD",x"9F",x"28",x"CD", -- 0x2B28
		x"DC",x"2C",x"CD",x"9A",x"26",x"21",x"11",x"2D", -- 0x2B30
		x"CD",x"3B",x"2C",x"CD",x"4D",x"2C",x"CD",x"E1", -- 0x2B38
		x"2C",x"3A",x"9D",x"F6",x"3D",x"20",x"DC",x"C3", -- 0x2B40
		x"59",x"2C",x"21",x"09",x"2D",x"CD",x"3B",x"2C", -- 0x2B48
		x"CD",x"CC",x"2C",x"CD",x"8A",x"2F",x"7D",x"17", -- 0x2B50
		x"9F",x"BC",x"28",x"14",x"7C",x"B7",x"F2",x"6D", -- 0x2B58
		x"2B",x"CD",x"4F",x"30",x"CD",x"E1",x"2C",x"21", -- 0x2B60
		x"13",x"2D",x"C3",x"5C",x"2C",x"C3",x"67",x"40", -- 0x2B68
		x"22",x"9D",x"F6",x"CD",x"3A",x"30",x"CD",x"4D", -- 0x2B70
		x"2C",x"CD",x"E1",x"2C",x"CD",x"8C",x"26",x"21", -- 0x2B78
		x"11",x"2D",x"CD",x"47",x"2C",x"F5",x"28",x"08", -- 0x2B80
		x"38",x"06",x"21",x"11",x"2D",x"CD",x"32",x"2C", -- 0x2B88
		x"CD",x"CC",x"2C",x"21",x"8C",x"2D",x"CD",x"88", -- 0x2B90
		x"2C",x"CD",x"6F",x"2C",x"21",x"6B",x"2D",x"CD", -- 0x2B98
		x"9A",x"2C",x"CD",x"DC",x"2C",x"CD",x"C7",x"2C", -- 0x2BA0
		x"CD",x"CC",x"2C",x"CD",x"8C",x"26",x"21",x"3E", -- 0x2BA8
		x"F8",x"CD",x"67",x"2C",x"CD",x"DC",x"2C",x"CD", -- 0x2BB0
		x"E1",x"2C",x"CD",x"9A",x"26",x"21",x"3E",x"F8", -- 0x2BB8
		x"CD",x"50",x"2C",x"CD",x"9F",x"28",x"F1",x"38", -- 0x2BC0
		x"08",x"28",x"06",x"21",x"2B",x"2D",x"CD",x"3B", -- 0x2BC8
		x"2C",x"3A",x"9D",x"F6",x"21",x"F6",x"F7",x"4E", -- 0x2BD0
		x"86",x"77",x"A9",x"F0",x"C3",x"67",x"40",x"CD", -- 0x2BD8
		x"71",x"2E",x"21",x"57",x"F8",x"28",x"2E",x"FC", -- 0x2BE0
		x"67",x"2C",x"21",x"3E",x"F8",x"11",x"57",x"F8", -- 0x2BE8
		x"CD",x"6A",x"2C",x"21",x"F9",x"2C",x"CD",x"50", -- 0x2BF0
		x"2C",x"21",x"F1",x"2C",x"CD",x"5C",x"2C",x"11", -- 0x2BF8
		x"45",x"F8",x"CD",x"2E",x"28",x"11",x"FE",x"F7", -- 0x2C00
		x"21",x"58",x"F8",x"06",x"07",x"CD",x"F7",x"2E", -- 0x2C08
		x"21",x"57",x"F8",x"36",x"00",x"CD",x"5C",x"2C", -- 0x2C10
		x"21",x"F6",x"F7",x"36",x"40",x"AF",x"32",x"FE", -- 0x2C18
		x"F7",x"C3",x"FA",x"26",x"11",x"01",x"2D",x"21", -- 0x2C20
		x"57",x"F8",x"18",x"3E",x"CD",x"50",x"2C",x"C3", -- 0x2C28
		x"9A",x"26",x"CD",x"50",x"2C",x"C3",x"8C",x"26", -- 0x2C30
		x"21",x"F6",x"F7",x"CD",x"50",x"2C",x"C3",x"E6", -- 0x2C38
		x"27",x"CD",x"50",x"2C",x"C3",x"9F",x"28",x"CD", -- 0x2C40
		x"50",x"2C",x"C3",x"5C",x"2F",x"21",x"F6",x"F7", -- 0x2C48
		x"11",x"47",x"F8",x"EB",x"CD",x"6A",x"2C",x"EB", -- 0x2C50
		x"C9",x"21",x"47",x"F8",x"11",x"F6",x"F7",x"18", -- 0x2C58
		x"F2",x"CD",x"CB",x"2F",x"21",x"57",x"F8",x"11", -- 0x2C60
		x"F6",x"F7",x"06",x"08",x"C3",x"F7",x"2E",x"E1", -- 0x2C68
		x"22",x"C5",x"F7",x"CD",x"DC",x"2C",x"CD",x"CC", -- 0x2C70
		x"2C",x"CD",x"59",x"2C",x"2A",x"C5",x"F7",x"E9", -- 0x2C78
		x"CD",x"8D",x"2E",x"21",x"8D",x"2E",x"E3",x"E9", -- 0x2C80
		x"22",x"C5",x"F7",x"CD",x"CC",x"2C",x"2A",x"C5", -- 0x2C88
		x"F7",x"CD",x"9A",x"2C",x"CD",x"DC",x"2C",x"C3", -- 0x2C90
		x"E6",x"27",x"22",x"C5",x"F7",x"CD",x"38",x"2C", -- 0x2C98
		x"2A",x"C5",x"F7",x"7E",x"F5",x"23",x"E5",x"21", -- 0x2CA0
		x"C5",x"F7",x"CD",x"67",x"2C",x"E1",x"CD",x"5C", -- 0x2CA8
		x"2C",x"F1",x"3D",x"C8",x"F5",x"E5",x"21",x"C5", -- 0x2CB0
		x"F7",x"CD",x"3B",x"2C",x"E1",x"CD",x"50",x"2C", -- 0x2CB8
		x"E5",x"CD",x"9A",x"26",x"E1",x"18",x"EA",x"21", -- 0x2CC0
		x"4E",x"F8",x"18",x"03",x"21",x"FD",x"F7",x"3E", -- 0x2CC8
		x"04",x"D1",x"46",x"2B",x"4E",x"2B",x"C5",x"3D", -- 0x2CD0
		x"20",x"F8",x"EB",x"E9",x"21",x"47",x"F8",x"18", -- 0x2CD8
		x"03",x"21",x"F6",x"F7",x"3E",x"04",x"D1",x"C1", -- 0x2CE0
		x"71",x"23",x"70",x"23",x"3D",x"20",x"F8",x"EB", -- 0x2CE8
		x"E9",x"00",x"14",x"38",x"98",x"20",x"42",x"08", -- 0x2CF0
		x"21",x"00",x"21",x"13",x"24",x"86",x"54",x"05", -- 0x2CF8
		x"19",x"00",x"40",x"64",x"96",x"51",x"37",x"23", -- 0x2D00
		x"58",x"40",x"43",x"42",x"94",x"48",x"19",x"03", -- 0x2D08
		x"24",x"40",x"50",x"00",x"00",x"00",x"00",x"00", -- 0x2D10
		x"00",x"00",x"00",x"41",x"10",x"00",x"00",x"00", -- 0x2D18
		x"00",x"00",x"00",x"40",x"25",x"00",x"00",x"00", -- 0x2D20
		x"00",x"00",x"00",x"41",x"31",x"62",x"27",x"76", -- 0x2D28
		x"60",x"16",x"84",x"40",x"86",x"85",x"88",x"96", -- 0x2D30
		x"38",x"06",x"50",x"41",x"23",x"02",x"58",x"50", -- 0x2D38
		x"92",x"99",x"40",x"41",x"15",x"70",x"79",x"63", -- 0x2D40
		x"26",x"79",x"49",x"40",x"26",x"79",x"49",x"19", -- 0x2D48
		x"24",x"31",x"12",x"41",x"17",x"32",x"05",x"08", -- 0x2D50
		x"07",x"56",x"89",x"40",x"52",x"35",x"98",x"77", -- 0x2D58
		x"55",x"98",x"30",x"40",x"15",x"91",x"54",x"94", -- 0x2D60
		x"30",x"91",x"90",x"04",x"41",x"10",x"00",x"00", -- 0x2D68
		x"00",x"00",x"00",x"00",x"43",x"15",x"93",x"74", -- 0x2D70
		x"15",x"23",x"60",x"31",x"44",x"27",x"09",x"31", -- 0x2D78
		x"69",x"40",x"85",x"16",x"44",x"44",x"97",x"63", -- 0x2D80
		x"35",x"57",x"40",x"58",x"03",x"42",x"18",x"31", -- 0x2D88
		x"23",x"60",x"15",x"92",x"75",x"43",x"83",x"14", -- 0x2D90
		x"06",x"72",x"12",x"93",x"71",x"44",x"51",x"78", -- 0x2D98
		x"09",x"19",x"91",x"51",x"62",x"04",x"C0",x"71", -- 0x2DA0
		x"43",x"33",x"82",x"15",x"32",x"26",x"41",x"62", -- 0x2DA8
		x"50",x"36",x"51",x"12",x"79",x"08",x"C2",x"13", -- 0x2DB0
		x"68",x"23",x"70",x"24",x"15",x"03",x"41",x"85", -- 0x2DB8
		x"16",x"73",x"19",x"87",x"23",x"89",x"05",x"41", -- 0x2DC0
		x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"C2", -- 0x2DC8
		x"13",x"21",x"04",x"78",x"35",x"01",x"56",x"42", -- 0x2DD0
		x"47",x"92",x"52",x"56",x"04",x"38",x"73",x"C2", -- 0x2DD8
		x"64",x"90",x"66",x"82",x"74",x"09",x"43",x"42", -- 0x2DE0
		x"29",x"41",x"57",x"50",x"17",x"23",x"23",x"08", -- 0x2DE8
		x"C0",x"69",x"21",x"56",x"92",x"29",x"18",x"09", -- 0x2DF0
		x"41",x"38",x"17",x"28",x"86",x"38",x"57",x"71", -- 0x2DF8
		x"C2",x"15",x"09",x"44",x"99",x"47",x"48",x"01", -- 0x2E00
		x"42",x"42",x"05",x"86",x"89",x"66",x"73",x"55", -- 0x2E08
		x"C2",x"76",x"70",x"58",x"59",x"68",x"32",x"91", -- 0x2E10
		x"42",x"81",x"60",x"52",x"49",x"27",x"55",x"13", -- 0x2E18
		x"C2",x"41",x"34",x"17",x"02",x"24",x"03",x"98", -- 0x2E20
		x"41",x"62",x"83",x"18",x"53",x"07",x"17",x"96", -- 0x2E28
		x"08",x"BF",x"52",x"08",x"69",x"39",x"04",x"00", -- 0x2E30
		x"00",x"3F",x"75",x"30",x"71",x"49",x"13",x"48", -- 0x2E38
		x"00",x"BF",x"90",x"81",x"34",x"32",x"24",x"70", -- 0x2E40
		x"50",x"40",x"11",x"11",x"07",x"94",x"18",x"40", -- 0x2E48
		x"29",x"C0",x"14",x"28",x"57",x"08",x"55",x"48", -- 0x2E50
		x"84",x"40",x"19",x"99",x"99",x"99",x"94",x"89", -- 0x2E58
		x"67",x"C0",x"33",x"33",x"33",x"33",x"33",x"31", -- 0x2E60
		x"60",x"41",x"10",x"00",x"00",x"00",x"00",x"00", -- 0x2E68
		x"00",x"3A",x"F6",x"F7",x"B7",x"C8",x"FE",x"2F", -- 0x2E70
		x"17",x"9F",x"C0",x"3C",x"C9",x"AF",x"32",x"F6", -- 0x2E78
		x"F7",x"C9",x"CD",x"A1",x"2E",x"F0",x"EF",x"FA", -- 0x2E80
		x"2B",x"32",x"CA",x"6D",x"40",x"21",x"F6",x"F7", -- 0x2E88
		x"7E",x"B7",x"C8",x"EE",x"80",x"77",x"C9",x"CD", -- 0x2E90
		x"A1",x"2E",x"6F",x"17",x"9F",x"67",x"C3",x"99", -- 0x2E98
		x"2F",x"EF",x"CA",x"6D",x"40",x"F2",x"71",x"2E", -- 0x2EA0
		x"2A",x"F8",x"F7",x"7C",x"B5",x"C8",x"7C",x"18", -- 0x2EA8
		x"C7",x"EB",x"2A",x"F8",x"F7",x"E3",x"E5",x"2A", -- 0x2EB0
		x"F6",x"F7",x"E3",x"E5",x"EB",x"C9",x"CD",x"DF", -- 0x2EB8
		x"2E",x"EB",x"22",x"F8",x"F7",x"60",x"69",x"22", -- 0x2EC0
		x"F6",x"F7",x"EB",x"C9",x"2A",x"F8",x"F7",x"EB", -- 0x2EC8
		x"2A",x"F6",x"F7",x"4D",x"44",x"C9",x"4E",x"23", -- 0x2ED0
		x"46",x"23",x"5E",x"23",x"56",x"23",x"C9",x"5E", -- 0x2ED8
		x"23",x"56",x"23",x"4E",x"23",x"46",x"23",x"C9", -- 0x2EE0
		x"11",x"F6",x"F7",x"06",x"04",x"18",x"08",x"11", -- 0x2EE8
		x"47",x"F8",x"EB",x"3A",x"63",x"F6",x"47",x"1A", -- 0x2EF0
		x"77",x"13",x"23",x"10",x"FA",x"C9",x"1A",x"77", -- 0x2EF8
		x"1B",x"2B",x"10",x"FA",x"C9",x"21",x"47",x"F8", -- 0x2F00
		x"11",x"F2",x"2E",x"18",x"06",x"21",x"47",x"F8", -- 0x2F08
		x"11",x"F3",x"2E",x"D5",x"11",x"F6",x"F7",x"3A", -- 0x2F10
		x"63",x"F6",x"FE",x"04",x"D0",x"11",x"F8",x"F7", -- 0x2F18
		x"C9",x"79",x"B7",x"CA",x"71",x"2E",x"21",x"77", -- 0x2F20
		x"2E",x"E5",x"CD",x"71",x"2E",x"79",x"C8",x"21", -- 0x2F28
		x"F6",x"F7",x"AE",x"79",x"F8",x"CD",x"3B",x"2F", -- 0x2F30
		x"1F",x"A9",x"C9",x"79",x"BE",x"C0",x"23",x"78", -- 0x2F38
		x"BE",x"C0",x"23",x"7B",x"BE",x"C0",x"23",x"7A", -- 0x2F40
		x"96",x"C0",x"E1",x"E1",x"C9",x"7A",x"AC",x"7C", -- 0x2F48
		x"FA",x"78",x"2E",x"BA",x"20",x"03",x"7D",x"93", -- 0x2F50
		x"C8",x"C3",x"79",x"2E",x"11",x"47",x"F8",x"1A", -- 0x2F58
		x"B7",x"CA",x"71",x"2E",x"21",x"77",x"2E",x"E5", -- 0x2F60
		x"CD",x"71",x"2E",x"1A",x"4F",x"C8",x"21",x"F6", -- 0x2F68
		x"F7",x"AE",x"79",x"F8",x"06",x"08",x"1A",x"96", -- 0x2F70
		x"20",x"06",x"13",x"23",x"10",x"F8",x"C1",x"C9", -- 0x2F78
		x"1F",x"A9",x"C9",x"CD",x"5C",x"2F",x"C2",x"77", -- 0x2F80
		x"2E",x"C9",x"EF",x"2A",x"F8",x"F7",x"F8",x"CA", -- 0x2F88
		x"6D",x"40",x"CD",x"5D",x"30",x"DA",x"67",x"40", -- 0x2F90
		x"EB",x"22",x"F8",x"F7",x"3E",x"02",x"32",x"63", -- 0x2F98
		x"F6",x"C9",x"01",x"C5",x"32",x"11",x"76",x"80", -- 0x2FA0
		x"CD",x"21",x"2F",x"C0",x"21",x"00",x"80",x"D1", -- 0x2FA8
		x"18",x"E7",x"EF",x"E0",x"FA",x"C8",x"2F",x"CA", -- 0x2FB0
		x"6D",x"40",x"CD",x"53",x"30",x"CD",x"52",x"37", -- 0x2FB8
		x"23",x"78",x"B7",x"1F",x"47",x"C3",x"41",x"27", -- 0x2FC0
		x"2A",x"F8",x"F7",x"7C",x"B7",x"F5",x"FC",x"21", -- 0x2FC8
		x"32",x"CD",x"53",x"30",x"EB",x"21",x"00",x"00", -- 0x2FD0
		x"22",x"F6",x"F7",x"22",x"F8",x"F7",x"7A",x"B3", -- 0x2FD8
		x"CA",x"A7",x"66",x"01",x"00",x"05",x"21",x"F7", -- 0x2FE0
		x"F7",x"E5",x"21",x"30",x"30",x"3E",x"FF",x"D5", -- 0x2FE8
		x"5E",x"23",x"56",x"23",x"E3",x"C5",x"44",x"4D", -- 0x2FF0
		x"19",x"3C",x"38",x"FA",x"60",x"69",x"C1",x"D1", -- 0x2FF8
		x"EB",x"0C",x"0D",x"20",x"0B",x"B7",x"28",x"1C", -- 0x3000
		x"F5",x"3E",x"40",x"80",x"32",x"F6",x"F7",x"F1", -- 0x3008
		x"0C",x"E3",x"F5",x"79",x"1F",x"30",x"08",x"F1", -- 0x3010
		x"87",x"87",x"87",x"87",x"77",x"18",x"04",x"F1", -- 0x3018
		x"B6",x"77",x"23",x"E3",x"7A",x"B3",x"28",x"02", -- 0x3020
		x"10",x"C3",x"E1",x"F1",x"F0",x"C3",x"8D",x"2E", -- 0x3028
		x"F0",x"D8",x"18",x"FC",x"9C",x"FF",x"F6",x"FF", -- 0x3030
		x"FF",x"FF",x"EF",x"D0",x"CA",x"6D",x"40",x"FC", -- 0x3038
		x"C8",x"2F",x"21",x"00",x"00",x"22",x"FA",x"F7", -- 0x3040
		x"22",x"FC",x"F7",x"7C",x"32",x"FE",x"F7",x"3E", -- 0x3048
		x"08",x"18",x"02",x"3E",x"04",x"C3",x"9E",x"2F", -- 0x3050
		x"EF",x"C8",x"C3",x"6D",x"40",x"21",x"BA",x"30", -- 0x3058
		x"E5",x"21",x"F6",x"F7",x"7E",x"E6",x"7F",x"FE", -- 0x3060
		x"46",x"D0",x"D6",x"41",x"30",x"06",x"B7",x"D1", -- 0x3068
		x"11",x"00",x"00",x"C9",x"3C",x"47",x"11",x"00", -- 0x3070
		x"00",x"4A",x"23",x"79",x"0C",x"1F",x"7E",x"38", -- 0x3078
		x"06",x"1F",x"1F",x"1F",x"1F",x"18",x"01",x"23", -- 0x3080
		x"E6",x"0F",x"22",x"F0",x"F7",x"62",x"6B",x"29", -- 0x3088
		x"D8",x"29",x"D8",x"19",x"D8",x"29",x"D8",x"5F", -- 0x3090
		x"16",x"00",x"19",x"D8",x"EB",x"2A",x"F0",x"F7", -- 0x3098
		x"10",x"D9",x"21",x"00",x"80",x"E7",x"3A",x"F6", -- 0x30A0
		x"F7",x"D8",x"28",x"0A",x"E1",x"B7",x"F0",x"EB", -- 0x30A8
		x"CD",x"21",x"32",x"EB",x"B7",x"C9",x"B7",x"F0", -- 0x30B0
		x"E1",x"C9",x"37",x"C9",x"0B",x"C9",x"EF",x"F8", -- 0x30B8
		x"CD",x"71",x"2E",x"F2",x"CF",x"30",x"CD",x"8D", -- 0x30C0
		x"2E",x"CD",x"CF",x"30",x"C3",x"86",x"2E",x"EF", -- 0x30C8
		x"F8",x"21",x"FE",x"F7",x"0E",x"0E",x"30",x"08", -- 0x30D0
		x"CA",x"6D",x"40",x"21",x"FA",x"F7",x"0E",x"06", -- 0x30D8
		x"3A",x"F6",x"F7",x"B7",x"FA",x"00",x"31",x"E6", -- 0x30E0
		x"7F",x"D6",x"41",x"DA",x"7D",x"2E",x"3C",x"91", -- 0x30E8
		x"D0",x"2F",x"3C",x"47",x"2B",x"7E",x"E6",x"F0", -- 0x30F0
		x"77",x"05",x"C8",x"AF",x"77",x"10",x"F5",x"C9", -- 0x30F8
		x"E6",x"7F",x"D6",x"41",x"30",x"06",x"21",x"FF", -- 0x3100
		x"FF",x"C3",x"99",x"2F",x"3C",x"91",x"D0",x"2F", -- 0x3108
		x"3C",x"47",x"1E",x"00",x"2B",x"7E",x"57",x"E6", -- 0x3110
		x"F0",x"77",x"BA",x"28",x"01",x"1C",x"05",x"28", -- 0x3118
		x"08",x"AF",x"77",x"BA",x"28",x"01",x"1C",x"10", -- 0x3120
		x"EB",x"1C",x"1D",x"C8",x"79",x"FE",x"06",x"01", -- 0x3128
		x"C1",x"10",x"11",x"00",x"00",x"CA",x"4E",x"32", -- 0x3130
		x"EB",x"22",x"4D",x"F8",x"22",x"4B",x"F8",x"22", -- 0x3138
		x"49",x"F8",x"60",x"69",x"22",x"47",x"F8",x"C3", -- 0x3140
		x"9A",x"26",x"E5",x"21",x"00",x"00",x"78",x"B1", -- 0x3148
		x"28",x"12",x"3E",x"10",x"29",x"DA",x"1D",x"60", -- 0x3150
		x"EB",x"29",x"EB",x"30",x"04",x"09",x"DA",x"1D", -- 0x3158
		x"60",x"3D",x"20",x"F0",x"EB",x"E1",x"C9",x"7C", -- 0x3160
		x"17",x"9F",x"47",x"CD",x"21",x"32",x"79",x"98", -- 0x3168
		x"18",x"03",x"7C",x"17",x"9F",x"47",x"E5",x"7A", -- 0x3170
		x"17",x"9F",x"19",x"88",x"0F",x"AC",x"F2",x"AF", -- 0x3178
		x"2F",x"C5",x"EB",x"CD",x"CB",x"2F",x"F1",x"E1", -- 0x3180
		x"CD",x"B1",x"2E",x"CD",x"CB",x"2F",x"C1",x"D1", -- 0x3188
		x"C3",x"4E",x"32",x"7C",x"B5",x"CA",x"99",x"2F", -- 0x3190
		x"E5",x"D5",x"CD",x"15",x"32",x"C5",x"44",x"4D", -- 0x3198
		x"21",x"00",x"00",x"3E",x"10",x"29",x"38",x"1F", -- 0x31A0
		x"EB",x"29",x"EB",x"30",x"03",x"09",x"38",x"17", -- 0x31A8
		x"3D",x"20",x"F2",x"C1",x"D1",x"7C",x"B7",x"FA", -- 0x31B0
		x"BF",x"31",x"D1",x"78",x"C3",x"1D",x"32",x"EE", -- 0x31B8
		x"80",x"B5",x"28",x"14",x"EB",x"18",x"02",x"C1", -- 0x31C0
		x"E1",x"CD",x"CB",x"2F",x"E1",x"CD",x"B1",x"2E", -- 0x31C8
		x"CD",x"CB",x"2F",x"C1",x"D1",x"C3",x"5C",x"32", -- 0x31D0
		x"78",x"B7",x"C1",x"FA",x"99",x"2F",x"D5",x"CD", -- 0x31D8
		x"CB",x"2F",x"D1",x"C3",x"8D",x"2E",x"7C",x"B5", -- 0x31E0
		x"CA",x"58",x"40",x"CD",x"15",x"32",x"C5",x"EB", -- 0x31E8
		x"CD",x"21",x"32",x"44",x"4D",x"21",x"00",x"00", -- 0x31F0
		x"3E",x"11",x"B7",x"18",x"09",x"E5",x"09",x"30", -- 0x31F8
		x"04",x"33",x"33",x"37",x"30",x"E1",x"CB",x"13", -- 0x3200
		x"CB",x"12",x"ED",x"6A",x"3D",x"20",x"EE",x"EB", -- 0x3208
		x"C1",x"D5",x"C3",x"B5",x"31",x"7C",x"AA",x"47", -- 0x3210
		x"CD",x"1C",x"32",x"EB",x"7C",x"B7",x"F2",x"99", -- 0x3218
		x"2F",x"AF",x"4F",x"95",x"6F",x"79",x"9C",x"67", -- 0x3220
		x"C3",x"99",x"2F",x"2A",x"F8",x"F7",x"CD",x"21", -- 0x3228
		x"32",x"7C",x"EE",x"80",x"B5",x"C0",x"AF",x"C3", -- 0x3230
		x"CC",x"2F",x"D5",x"CD",x"E6",x"31",x"AF",x"82", -- 0x3238
		x"1F",x"67",x"7B",x"1F",x"6F",x"CD",x"9C",x"2F", -- 0x3240
		x"F1",x"18",x"D2",x"CD",x"DF",x"2E",x"CD",x"80", -- 0x3248
		x"32",x"CD",x"42",x"30",x"C3",x"9A",x"26",x"CD", -- 0x3250
		x"8D",x"2E",x"18",x"F2",x"CD",x"80",x"32",x"CD", -- 0x3258
		x"42",x"30",x"C3",x"E6",x"27",x"C1",x"D1",x"2A", -- 0x3260
		x"F8",x"F7",x"EB",x"22",x"F8",x"F7",x"C5",x"2A", -- 0x3268
		x"F6",x"F7",x"E3",x"22",x"F6",x"F7",x"C1",x"CD", -- 0x3270
		x"80",x"32",x"CD",x"42",x"30",x"C3",x"9F",x"28", -- 0x3278
		x"EB",x"22",x"49",x"F8",x"60",x"69",x"22",x"47", -- 0x3280
		x"F8",x"21",x"00",x"00",x"22",x"4B",x"F8",x"22", -- 0x3288
		x"4D",x"F8",x"C9",x"3D",x"C9",x"2B",x"C9",x"E1", -- 0x3290
		x"C9",x"EB",x"01",x"FF",x"00",x"60",x"68",x"CD", -- 0x3298
		x"99",x"2F",x"EB",x"7E",x"FE",x"26",x"CA",x"B8", -- 0x32A0
		x"4E",x"FE",x"2D",x"F5",x"28",x"05",x"FE",x"2B", -- 0x32A8
		x"28",x"01",x"2B",x"D7",x"DA",x"86",x"33",x"FE", -- 0x32B0
		x"2E",x"CA",x"4F",x"33",x"FE",x"65",x"28",x"02", -- 0x32B8
		x"FE",x"45",x"20",x"1A",x"E5",x"D7",x"FE",x"6C", -- 0x32C0
		x"28",x"0A",x"FE",x"4C",x"28",x"06",x"FE",x"71", -- 0x32C8
		x"28",x"02",x"FE",x"51",x"E1",x"28",x"06",x"EF", -- 0x32D0
		x"30",x"1B",x"AF",x"18",x"19",x"7E",x"FE",x"25", -- 0x32D8
		x"CA",x"62",x"33",x"FE",x"23",x"CA",x"70",x"33", -- 0x32E0
		x"FE",x"21",x"CA",x"71",x"33",x"FE",x"64",x"28", -- 0x32E8
		x"04",x"FE",x"44",x"20",x"29",x"B7",x"CD",x"77", -- 0x32F0
		x"33",x"D7",x"D5",x"16",x"00",x"CD",x"47",x"4F", -- 0x32F8
		x"4A",x"D1",x"D7",x"30",x"13",x"7B",x"FE",x"0C", -- 0x3300
		x"30",x"0A",x"07",x"07",x"83",x"07",x"86",x"D6", -- 0x3308
		x"30",x"5F",x"18",x"EE",x"1E",x"80",x"18",x"EA", -- 0x3310
		x"0C",x"20",x"03",x"AF",x"93",x"5F",x"EF",x"FA", -- 0x3318
		x"34",x"33",x"3A",x"F6",x"F7",x"B7",x"28",x"0C", -- 0x3320
		x"7A",x"90",x"83",x"C6",x"40",x"32",x"F6",x"F7", -- 0x3328
		x"B7",x"FC",x"4C",x"33",x"F1",x"E5",x"CC",x"86", -- 0x3330
		x"2E",x"EF",x"30",x"0B",x"E1",x"E8",x"E5",x"21", -- 0x3338
		x"97",x"32",x"E5",x"CD",x"A2",x"2F",x"C9",x"CD", -- 0x3340
		x"3C",x"27",x"E1",x"C9",x"C3",x"67",x"40",x"EF", -- 0x3348
		x"0C",x"20",x"CB",x"30",x"0A",x"CD",x"77",x"33", -- 0x3350
		x"3A",x"F6",x"F7",x"B7",x"20",x"01",x"57",x"C3", -- 0x3358
		x"B3",x"32",x"D7",x"F1",x"E5",x"21",x"97",x"32", -- 0x3360
		x"E5",x"21",x"8A",x"2F",x"E5",x"F5",x"18",x"AE", -- 0x3368
		x"B7",x"CD",x"77",x"33",x"D7",x"18",x"A7",x"E5", -- 0x3370
		x"D5",x"C5",x"F5",x"CC",x"B2",x"2F",x"F1",x"C4", -- 0x3378
		x"3A",x"30",x"C1",x"D1",x"E1",x"C9",x"D6",x"30", -- 0x3380
		x"C2",x"93",x"33",x"B1",x"CA",x"93",x"33",x"A2", -- 0x3388
		x"CA",x"B3",x"32",x"14",x"7A",x"FE",x"07",x"20", -- 0x3390
		x"04",x"B7",x"CD",x"77",x"33",x"D5",x"78",x"81", -- 0x3398
		x"3C",x"47",x"C5",x"E5",x"7E",x"D6",x"30",x"F5", -- 0x33A0
		x"EF",x"F2",x"D1",x"33",x"2A",x"F8",x"F7",x"11", -- 0x33A8
		x"CD",x"0C",x"E7",x"30",x"19",x"54",x"5D",x"29", -- 0x33B0
		x"29",x"19",x"29",x"F1",x"4F",x"09",x"7C",x"B7", -- 0x33B8
		x"FA",x"CC",x"33",x"22",x"F8",x"F7",x"E1",x"C1", -- 0x33C0
		x"D1",x"C3",x"B3",x"32",x"79",x"F5",x"CD",x"C8", -- 0x33C8
		x"2F",x"F1",x"E1",x"C1",x"D1",x"20",x"0C",x"3A", -- 0x33D0
		x"F6",x"F7",x"B7",x"3E",x"00",x"20",x"04",x"57", -- 0x33D8
		x"C3",x"B3",x"32",x"D5",x"C5",x"E5",x"F5",x"21", -- 0x33E0
		x"F6",x"F7",x"36",x"01",x"7A",x"FE",x"10",x"38", -- 0x33E8
		x"03",x"F1",x"18",x"D2",x"3C",x"B7",x"1F",x"06", -- 0x33F0
		x"00",x"4F",x"09",x"F1",x"4F",x"7A",x"1F",x"79", -- 0x33F8
		x"30",x"04",x"87",x"87",x"87",x"87",x"B6",x"77", -- 0x3400
		x"18",x"BC",x"E5",x"21",x"D2",x"3F",x"CD",x"78", -- 0x3408
		x"66",x"E1",x"01",x"77",x"66",x"C5",x"CD",x"99", -- 0x3410
		x"2F",x"AF",x"32",x"9D",x"F6",x"21",x"C6",x"F7", -- 0x3418
		x"36",x"20",x"B6",x"18",x"1C",x"AF",x"CD",x"5F", -- 0x3420
		x"37",x"E6",x"08",x"28",x"02",x"36",x"2B",x"EB", -- 0x3428
		x"CD",x"A1",x"2E",x"EB",x"F2",x"41",x"34",x"36", -- 0x3430
		x"2D",x"C5",x"E5",x"CD",x"86",x"2E",x"E1",x"C1", -- 0x3438
		x"B4",x"23",x"36",x"30",x"3A",x"9D",x"F6",x"57", -- 0x3440
		x"17",x"3A",x"63",x"F6",x"DA",x"F7",x"34",x"CA", -- 0x3448
		x"EF",x"34",x"FE",x"04",x"D2",x"A1",x"34",x"01", -- 0x3450
		x"00",x"00",x"CD",x"DB",x"36",x"21",x"C6",x"F7", -- 0x3458
		x"46",x"0E",x"20",x"3A",x"9D",x"F6",x"5F",x"E6", -- 0x3460
		x"20",x"28",x"0C",x"78",x"B9",x"0E",x"2A",x"20", -- 0x3468
		x"06",x"7B",x"E6",x"04",x"20",x"01",x"41",x"71", -- 0x3470
		x"D7",x"28",x"14",x"FE",x"45",x"28",x"10",x"FE", -- 0x3478
		x"44",x"28",x"0C",x"FE",x"30",x"28",x"F0",x"FE", -- 0x3480
		x"2C",x"28",x"EC",x"FE",x"2E",x"20",x"03",x"2B", -- 0x3488
		x"36",x"30",x"7B",x"E6",x"10",x"28",x"03",x"2B", -- 0x3490
		x"36",x"24",x"7B",x"E6",x"04",x"C0",x"2B",x"70", -- 0x3498
		x"C9",x"E5",x"CD",x"52",x"37",x"50",x"14",x"01", -- 0x34A0
		x"00",x"03",x"3A",x"F6",x"F7",x"D6",x"3F",x"38", -- 0x34A8
		x"08",x"14",x"BA",x"30",x"04",x"3C",x"47",x"3E", -- 0x34B0
		x"02",x"D6",x"02",x"E1",x"F5",x"CD",x"8E",x"36", -- 0x34B8
		x"36",x"30",x"CC",x"E6",x"2E",x"CD",x"B3",x"36", -- 0x34C0
		x"2B",x"7E",x"FE",x"30",x"28",x"FA",x"FE",x"2E", -- 0x34C8
		x"C4",x"E6",x"2E",x"F1",x"28",x"1A",x"36",x"45", -- 0x34D0
		x"23",x"36",x"2B",x"F2",x"E2",x"34",x"36",x"2D", -- 0x34D8
		x"2F",x"3C",x"06",x"2F",x"04",x"D6",x"0A",x"30", -- 0x34E0
		x"FB",x"C6",x"3A",x"23",x"70",x"23",x"77",x"23", -- 0x34E8
		x"36",x"00",x"EB",x"21",x"C6",x"F7",x"C9",x"23", -- 0x34F0
		x"C5",x"FE",x"04",x"7A",x"D2",x"66",x"35",x"1F", -- 0x34F8
		x"DA",x"EF",x"35",x"01",x"03",x"06",x"CD",x"86", -- 0x3500
		x"36",x"D1",x"7A",x"D6",x"05",x"F4",x"66",x"36", -- 0x3508
		x"CD",x"DB",x"36",x"7B",x"B7",x"CC",x"95",x"32", -- 0x3510
		x"3D",x"F4",x"66",x"36",x"E5",x"CD",x"5D",x"34", -- 0x3518
		x"E1",x"28",x"02",x"70",x"23",x"36",x"00",x"21", -- 0x3520
		x"C5",x"F7",x"23",x"3A",x"BC",x"F6",x"95",x"92", -- 0x3528
		x"C8",x"7E",x"FE",x"20",x"28",x"F4",x"FE",x"2A", -- 0x3530
		x"28",x"F0",x"2B",x"E5",x"F5",x"01",x"3C",x"35", -- 0x3538
		x"C5",x"D7",x"FE",x"2D",x"C8",x"FE",x"2B",x"C8", -- 0x3540
		x"FE",x"24",x"C8",x"C1",x"FE",x"30",x"20",x"0F", -- 0x3548
		x"23",x"D7",x"30",x"0B",x"2B",x"18",x"02",x"2B", -- 0x3550
		x"77",x"F1",x"28",x"FB",x"C1",x"18",x"CC",x"F1", -- 0x3558
		x"28",x"FD",x"E1",x"36",x"25",x"C9",x"E5",x"1F", -- 0x3560
		x"DA",x"F5",x"35",x"CD",x"52",x"37",x"50",x"3A", -- 0x3568
		x"F6",x"F7",x"D6",x"4F",x"38",x"0B",x"E1",x"C1", -- 0x3570
		x"CD",x"25",x"34",x"21",x"C5",x"F7",x"36",x"25", -- 0x3578
		x"C9",x"CD",x"71",x"2E",x"C4",x"A2",x"37",x"E1", -- 0x3580
		x"C1",x"FA",x"A6",x"35",x"C5",x"5F",x"78",x"92", -- 0x3588
		x"93",x"F4",x"66",x"36",x"CD",x"7A",x"36",x"CD", -- 0x3590
		x"B3",x"36",x"B3",x"C4",x"74",x"36",x"B3",x"C4", -- 0x3598
		x"A0",x"36",x"D1",x"C3",x"13",x"35",x"5F",x"79", -- 0x35A0
		x"B7",x"C4",x"93",x"32",x"83",x"FA",x"B1",x"35", -- 0x35A8
		x"AF",x"C5",x"F5",x"FC",x"7B",x"37",x"C1",x"7B", -- 0x35B0
		x"90",x"C1",x"5F",x"82",x"78",x"FA",x"CB",x"35", -- 0x35B8
		x"92",x"93",x"F4",x"66",x"36",x"C5",x"CD",x"7A", -- 0x35C0
		x"36",x"18",x"11",x"CD",x"66",x"36",x"79",x"CD", -- 0x35C8
		x"A3",x"36",x"4F",x"AF",x"92",x"93",x"CD",x"66", -- 0x35D0
		x"36",x"C5",x"47",x"4F",x"CD",x"B3",x"36",x"C1", -- 0x35D8
		x"B1",x"20",x"03",x"2A",x"BC",x"F6",x"83",x"3D", -- 0x35E0
		x"F4",x"66",x"36",x"50",x"C3",x"1C",x"35",x"E5", -- 0x35E8
		x"D5",x"CD",x"C8",x"2F",x"D1",x"CD",x"52",x"37", -- 0x35F0
		x"58",x"CD",x"71",x"2E",x"F5",x"C4",x"A2",x"37", -- 0x35F8
		x"F1",x"E1",x"C1",x"F5",x"79",x"B7",x"F5",x"C4", -- 0x3600
		x"93",x"32",x"80",x"4F",x"7A",x"E6",x"04",x"FE", -- 0x3608
		x"01",x"9F",x"57",x"81",x"4F",x"93",x"F5",x"F2", -- 0x3610
		x"28",x"36",x"CD",x"7B",x"37",x"20",x"09",x"E5", -- 0x3618
		x"CD",x"DB",x"27",x"21",x"F6",x"F7",x"34",x"E1", -- 0x3620
		x"F1",x"C5",x"F5",x"FA",x"2F",x"36",x"AF",x"2F", -- 0x3628
		x"3C",x"80",x"3C",x"82",x"47",x"0E",x"00",x"CC", -- 0x3630
		x"8E",x"36",x"CD",x"B3",x"36",x"F1",x"F4",x"6E", -- 0x3638
		x"36",x"CD",x"A0",x"36",x"C1",x"F1",x"20",x"0C", -- 0x3640
		x"CD",x"95",x"32",x"7E",x"FE",x"2E",x"C4",x"E6", -- 0x3648
		x"2E",x"22",x"BC",x"F6",x"F1",x"3A",x"F6",x"F7", -- 0x3650
		x"28",x"03",x"83",x"90",x"92",x"C5",x"CD",x"D6", -- 0x3658
		x"34",x"EB",x"D1",x"C3",x"1C",x"35",x"B7",x"C8", -- 0x3660
		x"3D",x"36",x"30",x"23",x"18",x"F9",x"20",x"04", -- 0x3668
		x"C8",x"CD",x"A0",x"36",x"36",x"30",x"23",x"3D", -- 0x3670
		x"18",x"F6",x"7B",x"82",x"3C",x"47",x"3C",x"D6", -- 0x3678
		x"03",x"30",x"FC",x"C6",x"05",x"4F",x"3A",x"9D", -- 0x3680
		x"F6",x"E6",x"40",x"C0",x"4F",x"C9",x"05",x"F2", -- 0x3688
		x"A1",x"36",x"22",x"BC",x"F6",x"36",x"2E",x"23", -- 0x3690
		x"36",x"30",x"04",x"48",x"20",x"F9",x"23",x"C9", -- 0x3698
		x"05",x"20",x"08",x"36",x"2E",x"22",x"BC",x"F6", -- 0x36A0
		x"23",x"48",x"C9",x"0D",x"C0",x"36",x"2C",x"23", -- 0x36A8
		x"0E",x"03",x"C9",x"D5",x"E5",x"C5",x"CD",x"52", -- 0x36B0
		x"37",x"78",x"C1",x"E1",x"11",x"F7",x"F7",x"37", -- 0x36B8
		x"F5",x"CD",x"A0",x"36",x"1A",x"30",x"06",x"1F", -- 0x36C0
		x"1F",x"1F",x"1F",x"18",x"01",x"13",x"E6",x"0F", -- 0x36C8
		x"C6",x"30",x"77",x"23",x"F1",x"3D",x"3F",x"20", -- 0x36D0
		x"E7",x"18",x"2F",x"D5",x"11",x"10",x"37",x"3E", -- 0x36D8
		x"05",x"CD",x"A0",x"36",x"C5",x"F5",x"E5",x"EB", -- 0x36E0
		x"4E",x"23",x"46",x"C5",x"23",x"E3",x"EB",x"2A", -- 0x36E8
		x"F8",x"F7",x"06",x"2F",x"04",x"7D",x"93",x"6F", -- 0x36F0
		x"7C",x"9A",x"67",x"30",x"F7",x"19",x"22",x"F8", -- 0x36F8
		x"F7",x"D1",x"E1",x"70",x"23",x"F1",x"C1",x"3D", -- 0x3700
		x"20",x"D7",x"CD",x"A0",x"36",x"77",x"D1",x"C9", -- 0x3708
		x"10",x"27",x"E8",x"03",x"64",x"00",x"0A",x"00", -- 0x3710
		x"01",x"00",x"06",x"01",x"18",x"06",x"06",x"03", -- 0x3718
		x"18",x"02",x"06",x"04",x"C5",x"CD",x"39",x"54", -- 0x3720
		x"11",x"D6",x"F7",x"AF",x"12",x"C1",x"4F",x"C5", -- 0x3728
		x"1B",x"A7",x"7C",x"1F",x"67",x"7D",x"1F",x"6F", -- 0x3730
		x"79",x"1F",x"4F",x"10",x"F4",x"C1",x"C5",x"07", -- 0x3738
		x"10",x"FD",x"C6",x"30",x"FE",x"3A",x"38",x"02", -- 0x3740
		x"C6",x"07",x"12",x"C1",x"7D",x"B4",x"20",x"DF", -- 0x3748
		x"EB",x"C9",x"EF",x"21",x"FD",x"F7",x"06",x"0E", -- 0x3750
		x"D0",x"21",x"F9",x"F7",x"06",x"06",x"C9",x"32", -- 0x3758
		x"9D",x"F6",x"F5",x"C5",x"D5",x"CD",x"3A",x"30", -- 0x3760
		x"21",x"13",x"2D",x"3A",x"F6",x"F7",x"A7",x"CC", -- 0x3768
		x"5C",x"2C",x"D1",x"C1",x"F1",x"21",x"C6",x"F7", -- 0x3770
		x"36",x"20",x"C9",x"E5",x"D5",x"C5",x"F5",x"2F", -- 0x3778
		x"3C",x"5F",x"3E",x"01",x"CA",x"9C",x"37",x"CD", -- 0x3780
		x"52",x"37",x"E5",x"CD",x"DB",x"27",x"1D",x"20", -- 0x3788
		x"FA",x"E1",x"23",x"78",x"0F",x"47",x"CD",x"41", -- 0x3790
		x"27",x"CD",x"B4",x"37",x"C1",x"80",x"C1",x"D1", -- 0x3798
		x"E1",x"C9",x"C5",x"E5",x"CD",x"52",x"37",x"3A", -- 0x37A0
		x"F6",x"F7",x"D6",x"40",x"90",x"32",x"F6",x"F7", -- 0x37A8
		x"E1",x"C1",x"B7",x"C9",x"C5",x"CD",x"52",x"37", -- 0x37B0
		x"7E",x"E6",x"0F",x"20",x"08",x"05",x"7E",x"B7", -- 0x37B8
		x"20",x"03",x"2B",x"10",x"F3",x"78",x"C1",x"C9", -- 0x37C0
		x"CD",x"80",x"32",x"CD",x"42",x"30",x"CD",x"C7", -- 0x37C8
		x"2C",x"CD",x"6F",x"2C",x"CD",x"DC",x"2C",x"3A", -- 0x37D0
		x"47",x"F8",x"B7",x"CA",x"43",x"38",x"67",x"3A", -- 0x37D8
		x"F6",x"F7",x"B7",x"CA",x"4D",x"38",x"CD",x"CC", -- 0x37E0
		x"2C",x"CD",x"1A",x"39",x"38",x"3C",x"EB",x"22", -- 0x37E8
		x"9F",x"F6",x"CD",x"4F",x"30",x"CD",x"DC",x"2C", -- 0x37F0
		x"CD",x"1A",x"39",x"CD",x"4F",x"30",x"2A",x"9F", -- 0x37F8
		x"F6",x"D2",x"5A",x"38",x"3A",x"47",x"F8",x"F5", -- 0x3800
		x"E5",x"CD",x"59",x"2C",x"21",x"C5",x"F7",x"CD", -- 0x3808
		x"67",x"2C",x"21",x"1B",x"2D",x"CD",x"5C",x"2C", -- 0x3810
		x"E1",x"7C",x"B7",x"F5",x"F2",x"26",x"38",x"AF", -- 0x3818
		x"4F",x"95",x"6F",x"79",x"9C",x"67",x"E5",x"C3", -- 0x3820
		x"94",x"38",x"CD",x"4F",x"30",x"CD",x"59",x"2C", -- 0x3828
		x"CD",x"6F",x"2C",x"CD",x"72",x"2A",x"CD",x"DC", -- 0x3830
		x"2C",x"CD",x"E6",x"27",x"C3",x"4A",x"2B",x"7C", -- 0x3838
		x"B5",x"20",x"06",x"21",x"01",x"00",x"C3",x"57", -- 0x3840
		x"38",x"7A",x"B3",x"20",x"0D",x"7C",x"17",x"30", -- 0x3848
		x"03",x"C3",x"58",x"40",x"21",x"00",x"00",x"C3", -- 0x3850
		x"99",x"2F",x"22",x"9F",x"F6",x"D5",x"7C",x"B7", -- 0x3858
		x"F5",x"FC",x"21",x"32",x"44",x"4D",x"21",x"01", -- 0x3860
		x"00",x"B7",x"78",x"1F",x"47",x"79",x"1F",x"4F", -- 0x3868
		x"30",x"05",x"CD",x"0D",x"39",x"20",x"4C",x"78", -- 0x3870
		x"B1",x"28",x"63",x"E5",x"62",x"6B",x"CD",x"0D", -- 0x3878
		x"39",x"EB",x"E1",x"28",x"E4",x"C5",x"E5",x"21", -- 0x3880
		x"C5",x"F7",x"CD",x"67",x"2C",x"E1",x"CD",x"CB", -- 0x3888
		x"2F",x"CD",x"42",x"30",x"C1",x"78",x"B7",x"1F", -- 0x3890
		x"47",x"79",x"1F",x"4F",x"30",x"08",x"C5",x"21", -- 0x3898
		x"C5",x"F7",x"CD",x"3B",x"2C",x"C1",x"78",x"B1", -- 0x38A0
		x"28",x"34",x"C5",x"CD",x"CC",x"2C",x"21",x"C5", -- 0x38A8
		x"F7",x"E5",x"CD",x"5C",x"2C",x"E1",x"E5",x"CD", -- 0x38B0
		x"3B",x"2C",x"E1",x"CD",x"67",x"2C",x"CD",x"E1", -- 0x38B8
		x"2C",x"18",x"D1",x"C5",x"D5",x"CD",x"3A",x"30", -- 0x38C0
		x"CD",x"4D",x"2C",x"E1",x"CD",x"CB",x"2F",x"CD", -- 0x38C8
		x"42",x"30",x"21",x"C5",x"F7",x"CD",x"67",x"2C", -- 0x38D0
		x"CD",x"59",x"2C",x"C1",x"18",x"C8",x"F1",x"C1", -- 0x38D8
		x"F0",x"3A",x"63",x"F6",x"FE",x"02",x"20",x"08", -- 0x38E0
		x"C5",x"CD",x"CB",x"2F",x"CD",x"42",x"30",x"C1", -- 0x38E8
		x"3A",x"F6",x"F7",x"B7",x"20",x"0B",x"2A",x"9F", -- 0x38F0
		x"F6",x"B4",x"F0",x"7D",x"0F",x"A0",x"C3",x"67", -- 0x38F8
		x"40",x"CD",x"4D",x"2C",x"21",x"1B",x"2D",x"CD", -- 0x3900
		x"5C",x"2C",x"C3",x"9F",x"28",x"C5",x"D5",x"CD", -- 0x3908
		x"93",x"31",x"3A",x"63",x"F6",x"FE",x"02",x"D1", -- 0x3910
		x"C1",x"C9",x"CD",x"59",x"2C",x"CD",x"C7",x"2C", -- 0x3918
		x"CD",x"CF",x"30",x"CD",x"DC",x"2C",x"CD",x"5C", -- 0x3920
		x"2F",x"37",x"C0",x"C3",x"5D",x"30",x"EA",x"63", -- 0x3928
		x"24",x"45",x"27",x"65",x"5B",x"48",x"6C",x"4B", -- 0x3930
		x"9F",x"5E",x"9F",x"4B",x"80",x"48",x"E8",x"47", -- 0x3938
		x"9E",x"47",x"E5",x"49",x"C9",x"63",x"B2",x"47", -- 0x3940
		x"21",x"48",x"5D",x"48",x"E3",x"63",x"24",x"4A", -- 0x3948
		x"AF",x"64",x"2E",x"52",x"86",x"62",x"E4",x"48", -- 0x3950
		x"1C",x"40",x"1D",x"50",x"23",x"54",x"24",x"64", -- 0x3958
		x"B7",x"6F",x"3F",x"70",x"16",x"40",x"1D",x"4A", -- 0x3960
		x"29",x"52",x"C3",x"00",x"C9",x"51",x"5D",x"48", -- 0x3968
		x"38",x"64",x"39",x"64",x"3E",x"64",x"77",x"64", -- 0x3970
		x"AA",x"49",x"5D",x"49",x"E2",x"53",x"B5",x"49", -- 0x3978
		x"68",x"54",x"18",x"47",x"1B",x"47",x"1E",x"47", -- 0x3980
		x"21",x"47",x"0E",x"4B",x"B7",x"6A",x"52",x"7C", -- 0x3988
		x"5B",x"77",x"58",x"77",x"14",x"6C",x"5D",x"6B", -- 0x3990
		x"5E",x"6B",x"2F",x"6C",x"48",x"7C",x"4D",x"7C", -- 0x3998
		x"A3",x"6B",x"2A",x"6C",x"11",x"5B",x"80",x"79", -- 0x39A0
		x"6E",x"5D",x"C5",x"59",x"C0",x"00",x"E5",x"73", -- 0x39A8
		x"EA",x"57",x"E5",x"57",x"CA",x"73",x"CC",x"79", -- 0x39B0
		x"E2",x"7B",x"48",x"7A",x"37",x"7B",x"5A",x"7B", -- 0x39B8
		x"A8",x"55",x"11",x"79",x"6C",x"78",x"4B",x"7E", -- 0x39C0
		x"B7",x"73",x"C6",x"6E",x"92",x"6E",x"16",x"7C", -- 0x39C8
		x"1B",x"7C",x"20",x"7C",x"25",x"7C",x"2A",x"7C", -- 0x39D0
		x"2F",x"7C",x"34",x"7C",x"66",x"77",x"61",x"68", -- 0x39D8
		x"91",x"68",x"9A",x"68",x"97",x"2E",x"CF",x"30", -- 0x39E0
		x"82",x"2E",x"FF",x"2A",x"DF",x"2B",x"AC",x"29", -- 0x39E8
		x"72",x"2A",x"4A",x"2B",x"93",x"29",x"FB",x"29", -- 0x39F0
		x"14",x"2A",x"F2",x"69",x"01",x"40",x"CC",x"4F", -- 0x39F8
		x"FF",x"67",x"04",x"66",x"BB",x"68",x"0B",x"68", -- 0x3A00
		x"1B",x"68",x"1C",x"54",x"F5",x"7B",x"48",x"68", -- 0x3A08
		x"F5",x"65",x"FA",x"65",x"C7",x"4F",x"FF",x"65", -- 0x3A10
		x"8A",x"2F",x"B2",x"2F",x"3A",x"30",x"BE",x"30", -- 0x3A18
		x"40",x"79",x"4C",x"79",x"5A",x"79",x"69",x"79", -- 0x3A20
		x"39",x"7C",x"39",x"6D",x"66",x"7C",x"6B",x"7C", -- 0x3A28
		x"70",x"7C",x"25",x"6D",x"03",x"6D",x"14",x"6D", -- 0x3A30
		x"57",x"7C",x"5C",x"7C",x"61",x"7C",x"72",x"3A", -- 0x3A38
		x"88",x"3A",x"9F",x"3A",x"F3",x"3A",x"2E",x"3B", -- 0x3A40
		x"4F",x"3B",x"69",x"3B",x"7B",x"3B",x"80",x"3B", -- 0x3A48
		x"9F",x"3B",x"A0",x"3B",x"A8",x"3B",x"E8",x"3B", -- 0x3A50
		x"09",x"3C",x"18",x"3C",x"2B",x"3C",x"5D",x"3C", -- 0x3A58
		x"5E",x"3C",x"8E",x"3C",x"DB",x"3C",x"F6",x"3C", -- 0x3A60
		x"FF",x"3C",x"16",x"3D",x"20",x"3D",x"24",x"3D", -- 0x3A68
		x"25",x"3D",x"55",x"54",x"CF",x"A9",x"4E",x"C4", -- 0x3A70
		x"F6",x"42",x"D3",x"06",x"54",x"CE",x"0E",x"53", -- 0x3A78
		x"C3",x"15",x"54",x"54",x"52",x"A4",x"E9",x"00", -- 0x3A80
		x"41",x"53",x"C5",x"C9",x"53",x"41",x"56",x"C5", -- 0x3A88
		x"D0",x"4C",x"4F",x"41",x"C4",x"CF",x"45",x"45", -- 0x3A90
		x"D0",x"C0",x"49",x"4E",x"A4",x"1D",x"00",x"41", -- 0x3A98
		x"4C",x"CC",x"CA",x"4C",x"4F",x"53",x"C5",x"B4", -- 0x3AA0
		x"4F",x"50",x"D9",x"D6",x"4F",x"4E",x"D4",x"99", -- 0x3AA8
		x"4C",x"45",x"41",x"D2",x"92",x"4C",x"4F",x"41", -- 0x3AB0
		x"C4",x"9B",x"53",x"41",x"56",x"C5",x"9A",x"53", -- 0x3AB8
		x"52",x"4C",x"49",x"CE",x"E8",x"49",x"4E",x"D4", -- 0x3AC0
		x"1E",x"53",x"4E",x"C7",x"1F",x"44",x"42",x"CC", -- 0x3AC8
		x"20",x"56",x"C9",x"28",x"56",x"D3",x"29",x"56", -- 0x3AD0
		x"C4",x"2A",x"4F",x"D3",x"0C",x"48",x"52",x"A4", -- 0x3AD8
		x"16",x"49",x"52",x"43",x"4C",x"C5",x"BC",x"4F", -- 0x3AE0
		x"4C",x"4F",x"D2",x"BD",x"4C",x"D3",x"9F",x"4D", -- 0x3AE8
		x"C4",x"D7",x"00",x"45",x"4C",x"45",x"54",x"C5", -- 0x3AF0
		x"A8",x"41",x"54",x"C1",x"84",x"49",x"CD",x"86", -- 0x3AF8
		x"45",x"46",x"53",x"54",x"D2",x"AB",x"45",x"46", -- 0x3B00
		x"49",x"4E",x"D4",x"AC",x"45",x"46",x"53",x"4E", -- 0x3B08
		x"C7",x"AD",x"45",x"46",x"44",x"42",x"CC",x"AE", -- 0x3B10
		x"53",x"4B",x"4F",x"A4",x"D1",x"45",x"C6",x"97", -- 0x3B18
		x"53",x"4B",x"49",x"A4",x"EA",x"53",x"4B",x"C6", -- 0x3B20
		x"26",x"52",x"41",x"D7",x"BE",x"00",x"4C",x"53", -- 0x3B28
		x"C5",x"A1",x"4E",x"C4",x"81",x"52",x"41",x"53", -- 0x3B30
		x"C5",x"A5",x"52",x"52",x"4F",x"D2",x"A6",x"52", -- 0x3B38
		x"CC",x"E1",x"52",x"D2",x"E2",x"58",x"D0",x"0B", -- 0x3B40
		x"4F",x"C6",x"2B",x"51",x"D6",x"F9",x"00",x"4F", -- 0x3B48
		x"D2",x"82",x"49",x"45",x"4C",x"C4",x"B1",x"49", -- 0x3B50
		x"4C",x"45",x"D3",x"B7",x"CE",x"DE",x"52",x"C5", -- 0x3B58
		x"0F",x"49",x"D8",x"21",x"50",x"4F",x"D3",x"27", -- 0x3B60
		x"00",x"4F",x"54",x"CF",x"89",x"4F",x"20",x"54", -- 0x3B68
		x"CF",x"89",x"4F",x"53",x"55",x"C2",x"8D",x"45", -- 0x3B70
		x"D4",x"B2",x"00",x"45",x"58",x"A4",x"1B",x"00", -- 0x3B78
		x"4E",x"50",x"55",x"D4",x"85",x"C6",x"8B",x"4E", -- 0x3B80
		x"53",x"54",x"D2",x"E5",x"4E",x"D4",x"05",x"4E", -- 0x3B88
		x"D0",x"10",x"4D",x"D0",x"FA",x"4E",x"4B",x"45", -- 0x3B90
		x"59",x"A4",x"EC",x"50",x"CC",x"D5",x"00",x"00", -- 0x3B98
		x"49",x"4C",x"CC",x"D4",x"45",x"D9",x"CC",x"00", -- 0x3BA0
		x"50",x"52",x"49",x"4E",x"D4",x"9D",x"4C",x"49", -- 0x3BA8
		x"53",x"D4",x"9E",x"50",x"4F",x"D3",x"1C",x"45", -- 0x3BB0
		x"D4",x"88",x"4F",x"43",x"41",x"54",x"C5",x"D8", -- 0x3BB8
		x"49",x"4E",x"C5",x"AF",x"4F",x"41",x"C4",x"B5", -- 0x3BC0
		x"53",x"45",x"D4",x"B8",x"49",x"53",x"D4",x"93", -- 0x3BC8
		x"46",x"49",x"4C",x"45",x"D3",x"BB",x"4F",x"C7", -- 0x3BD0
		x"0A",x"4F",x"C3",x"2C",x"45",x"CE",x"12",x"45", -- 0x3BD8
		x"46",x"54",x"A4",x"01",x"4F",x"C6",x"2D",x"00", -- 0x3BE0
		x"4F",x"54",x"4F",x"D2",x"CE",x"45",x"52",x"47", -- 0x3BE8
		x"C5",x"B6",x"4F",x"C4",x"FB",x"4B",x"49",x"A4", -- 0x3BF0
		x"2E",x"4B",x"53",x"A4",x"2F",x"4B",x"44",x"A4", -- 0x3BF8
		x"30",x"49",x"44",x"A4",x"03",x"41",x"D8",x"CD", -- 0x3C00
		x"00",x"45",x"58",x"D4",x"83",x"41",x"4D",x"C5", -- 0x3C08
		x"D3",x"45",x"D7",x"94",x"4F",x"D4",x"E0",x"00", -- 0x3C10
		x"50",x"45",x"CE",x"B0",x"55",x"D4",x"9C",x"CE", -- 0x3C18
		x"95",x"D2",x"F7",x"43",x"54",x"A4",x"1A",x"46", -- 0x3C20
		x"C6",x"EB",x"00",x"52",x"49",x"4E",x"D4",x"91", -- 0x3C28
		x"55",x"D4",x"B3",x"4F",x"4B",x"C5",x"98",x"4F", -- 0x3C30
		x"D3",x"11",x"45",x"45",x"CB",x"17",x"53",x"45", -- 0x3C38
		x"D4",x"C2",x"52",x"45",x"53",x"45",x"D4",x"C3", -- 0x3C40
		x"4F",x"49",x"4E",x"D4",x"ED",x"41",x"49",x"4E", -- 0x3C48
		x"D4",x"BF",x"44",x"CC",x"24",x"41",x"C4",x"25", -- 0x3C50
		x"4C",x"41",x"D9",x"C1",x"00",x"00",x"45",x"54", -- 0x3C58
		x"55",x"52",x"CE",x"8E",x"45",x"41",x"C4",x"87", -- 0x3C60
		x"55",x"CE",x"8A",x"45",x"53",x"54",x"4F",x"52", -- 0x3C68
		x"C5",x"8C",x"45",x"CD",x"8F",x"45",x"53",x"55", -- 0x3C70
		x"4D",x"C5",x"A7",x"53",x"45",x"D4",x"B9",x"49", -- 0x3C78
		x"47",x"48",x"54",x"A4",x"02",x"4E",x"C4",x"08", -- 0x3C80
		x"45",x"4E",x"55",x"CD",x"AA",x"00",x"43",x"52", -- 0x3C88
		x"45",x"45",x"CE",x"C5",x"50",x"52",x"49",x"54", -- 0x3C90
		x"C5",x"C7",x"54",x"4F",x"D0",x"90",x"57",x"41", -- 0x3C98
		x"D0",x"A4",x"45",x"D4",x"D2",x"41",x"56",x"C5", -- 0x3CA0
		x"BA",x"50",x"43",x"A8",x"DF",x"54",x"45",x"D0", -- 0x3CA8
		x"DC",x"47",x"CE",x"04",x"51",x"D2",x"07",x"49", -- 0x3CB0
		x"CE",x"09",x"54",x"52",x"A4",x"13",x"54",x"52", -- 0x3CB8
		x"49",x"4E",x"47",x"A4",x"E3",x"50",x"41",x"43", -- 0x3CC0
		x"45",x"A4",x"19",x"4F",x"55",x"4E",x"C4",x"C4", -- 0x3CC8
		x"54",x"49",x"43",x"CB",x"22",x"54",x"52",x"49", -- 0x3CD0
		x"C7",x"23",x"00",x"48",x"45",x"CE",x"DA",x"52", -- 0x3CD8
		x"4F",x"CE",x"A2",x"52",x"4F",x"46",x"C6",x"A3", -- 0x3CE0
		x"41",x"42",x"A8",x"DB",x"CF",x"D9",x"49",x"4D", -- 0x3CE8
		x"C5",x"CB",x"41",x"CE",x"0D",x"00",x"53",x"49", -- 0x3CF0
		x"4E",x"C7",x"E4",x"53",x"D2",x"DD",x"00",x"41", -- 0x3CF8
		x"CC",x"14",x"41",x"52",x"50",x"54",x"D2",x"E7", -- 0x3D00
		x"44",x"D0",x"C8",x"50",x"4F",x"4B",x"C5",x"C6", -- 0x3D08
		x"50",x"45",x"45",x"CB",x"18",x"00",x"49",x"44", -- 0x3D10
		x"54",x"C8",x"A0",x"41",x"49",x"D4",x"96",x"00", -- 0x3D18
		x"4F",x"D2",x"F8",x"00",x"00",x"00",x"AB",x"F1", -- 0x3D20
		x"AD",x"F2",x"AA",x"F3",x"AF",x"F4",x"DE",x"F5", -- 0x3D28
		x"DC",x"FC",x"A7",x"E6",x"BE",x"EE",x"BD",x"EF", -- 0x3D30
		x"BC",x"F0",x"00",x"79",x"79",x"7C",x"7C",x"7F", -- 0x3D38
		x"50",x"46",x"3C",x"32",x"28",x"7A",x"7B",x"3A", -- 0x3D40
		x"30",x"00",x"00",x"8A",x"2F",x"58",x"30",x"B2", -- 0x3D48
		x"2F",x"9A",x"26",x"8C",x"26",x"E6",x"27",x"9F", -- 0x3D50
		x"28",x"D7",x"37",x"83",x"2F",x"4E",x"32",x"57", -- 0x3D58
		x"32",x"5C",x"32",x"67",x"32",x"C8",x"37",x"21", -- 0x3D60
		x"2F",x"72",x"31",x"67",x"31",x"93",x"31",x"B8", -- 0x3D68
		x"4D",x"3F",x"38",x"4D",x"2F",x"00",x"4E",x"45", -- 0x3D70
		x"58",x"54",x"20",x"77",x"69",x"74",x"68",x"6F", -- 0x3D78
		x"75",x"74",x"20",x"46",x"4F",x"52",x"00",x"53", -- 0x3D80
		x"79",x"6E",x"74",x"61",x"78",x"20",x"65",x"72", -- 0x3D88
		x"72",x"6F",x"72",x"00",x"52",x"45",x"54",x"55", -- 0x3D90
		x"52",x"4E",x"20",x"77",x"69",x"74",x"68",x"6F", -- 0x3D98
		x"75",x"74",x"20",x"47",x"4F",x"53",x"55",x"42", -- 0x3DA0
		x"00",x"4F",x"75",x"74",x"20",x"6F",x"66",x"20", -- 0x3DA8
		x"44",x"41",x"54",x"41",x"00",x"49",x"6C",x"6C", -- 0x3DB0
		x"65",x"67",x"61",x"6C",x"20",x"66",x"75",x"6E", -- 0x3DB8
		x"63",x"74",x"69",x"6F",x"6E",x"20",x"63",x"61", -- 0x3DC0
		x"6C",x"6C",x"00",x"4F",x"76",x"65",x"72",x"66", -- 0x3DC8
		x"6C",x"6F",x"77",x"00",x"4F",x"75",x"74",x"20", -- 0x3DD0
		x"6F",x"66",x"20",x"6D",x"65",x"6D",x"6F",x"72", -- 0x3DD8
		x"79",x"00",x"55",x"6E",x"64",x"65",x"66",x"69", -- 0x3DE0
		x"6E",x"65",x"64",x"20",x"6C",x"69",x"6E",x"65", -- 0x3DE8
		x"20",x"6E",x"75",x"6D",x"62",x"65",x"72",x"00", -- 0x3DF0
		x"53",x"75",x"62",x"73",x"63",x"72",x"69",x"70", -- 0x3DF8
		x"74",x"20",x"6F",x"75",x"74",x"20",x"6F",x"66", -- 0x3E00
		x"20",x"72",x"61",x"6E",x"67",x"65",x"00",x"52", -- 0x3E08
		x"65",x"64",x"69",x"6D",x"65",x"6E",x"73",x"69", -- 0x3E10
		x"6F",x"6E",x"65",x"64",x"20",x"61",x"72",x"72", -- 0x3E18
		x"61",x"79",x"00",x"44",x"69",x"76",x"69",x"73", -- 0x3E20
		x"69",x"6F",x"6E",x"20",x"62",x"79",x"20",x"7A", -- 0x3E28
		x"65",x"72",x"6F",x"00",x"49",x"6C",x"6C",x"65", -- 0x3E30
		x"67",x"61",x"6C",x"20",x"64",x"69",x"72",x"65", -- 0x3E38
		x"63",x"74",x"00",x"54",x"79",x"70",x"65",x"20", -- 0x3E40
		x"6D",x"69",x"73",x"6D",x"61",x"74",x"63",x"68", -- 0x3E48
		x"00",x"4F",x"75",x"74",x"20",x"6F",x"66",x"20", -- 0x3E50
		x"73",x"74",x"72",x"69",x"6E",x"67",x"20",x"73", -- 0x3E58
		x"70",x"61",x"63",x"65",x"00",x"53",x"74",x"72", -- 0x3E60
		x"69",x"6E",x"67",x"20",x"74",x"6F",x"6F",x"20", -- 0x3E68
		x"6C",x"6F",x"6E",x"67",x"00",x"53",x"74",x"72", -- 0x3E70
		x"69",x"6E",x"67",x"20",x"66",x"6F",x"72",x"6D", -- 0x3E78
		x"75",x"6C",x"61",x"20",x"74",x"6F",x"6F",x"20", -- 0x3E80
		x"63",x"6F",x"6D",x"70",x"6C",x"65",x"78",x"00", -- 0x3E88
		x"43",x"61",x"6E",x"27",x"74",x"20",x"43",x"4F", -- 0x3E90
		x"4E",x"54",x"49",x"4E",x"55",x"45",x"00",x"55", -- 0x3E98
		x"6E",x"64",x"65",x"66",x"69",x"6E",x"65",x"64", -- 0x3EA0
		x"20",x"75",x"73",x"65",x"72",x"20",x"66",x"75", -- 0x3EA8
		x"6E",x"63",x"74",x"69",x"6F",x"6E",x"00",x"44", -- 0x3EB0
		x"65",x"76",x"69",x"63",x"65",x"20",x"49",x"2F", -- 0x3EB8
		x"4F",x"20",x"65",x"72",x"72",x"6F",x"72",x"00", -- 0x3EC0
		x"56",x"65",x"72",x"69",x"66",x"79",x"20",x"65", -- 0x3EC8
		x"72",x"72",x"6F",x"72",x"00",x"4E",x"6F",x"20", -- 0x3ED0
		x"52",x"45",x"53",x"55",x"4D",x"45",x"00",x"52", -- 0x3ED8
		x"45",x"53",x"55",x"4D",x"45",x"20",x"77",x"69", -- 0x3EE0
		x"74",x"68",x"6F",x"75",x"74",x"20",x"65",x"72", -- 0x3EE8
		x"72",x"6F",x"72",x"00",x"55",x"6E",x"70",x"72", -- 0x3EF0
		x"69",x"6E",x"74",x"61",x"62",x"6C",x"65",x"20", -- 0x3EF8
		x"65",x"72",x"72",x"6F",x"72",x"00",x"4D",x"69", -- 0x3F00
		x"73",x"73",x"69",x"6E",x"67",x"20",x"6F",x"70", -- 0x3F08
		x"65",x"72",x"61",x"6E",x"64",x"00",x"4C",x"69", -- 0x3F10
		x"6E",x"65",x"20",x"62",x"75",x"66",x"66",x"65", -- 0x3F18
		x"72",x"20",x"6F",x"76",x"65",x"72",x"66",x"6C", -- 0x3F20
		x"6F",x"77",x"00",x"46",x"49",x"45",x"4C",x"44", -- 0x3F28
		x"20",x"6F",x"76",x"65",x"72",x"66",x"6C",x"6F", -- 0x3F30
		x"77",x"00",x"49",x"6E",x"74",x"65",x"72",x"6E", -- 0x3F38
		x"61",x"6C",x"20",x"65",x"72",x"72",x"6F",x"72", -- 0x3F40
		x"00",x"42",x"61",x"64",x"20",x"66",x"69",x"6C", -- 0x3F48
		x"65",x"20",x"6E",x"75",x"6D",x"62",x"65",x"72", -- 0x3F50
		x"00",x"46",x"69",x"6C",x"65",x"20",x"6E",x"6F", -- 0x3F58
		x"74",x"20",x"66",x"6F",x"75",x"6E",x"64",x"00", -- 0x3F60
		x"46",x"69",x"6C",x"65",x"20",x"61",x"6C",x"72", -- 0x3F68
		x"65",x"61",x"64",x"79",x"20",x"6F",x"70",x"65", -- 0x3F70
		x"6E",x"00",x"49",x"6E",x"70",x"75",x"74",x"20", -- 0x3F78
		x"70",x"61",x"73",x"74",x"20",x"65",x"6E",x"64", -- 0x3F80
		x"00",x"42",x"61",x"64",x"20",x"66",x"69",x"6C", -- 0x3F88
		x"65",x"20",x"6E",x"61",x"6D",x"65",x"00",x"44", -- 0x3F90
		x"69",x"72",x"65",x"63",x"74",x"20",x"73",x"74", -- 0x3F98
		x"61",x"74",x"65",x"6D",x"65",x"6E",x"74",x"20", -- 0x3FA0
		x"69",x"6E",x"20",x"66",x"69",x"6C",x"65",x"00", -- 0x3FA8
		x"53",x"65",x"71",x"75",x"65",x"6E",x"74",x"69", -- 0x3FB0
		x"61",x"6C",x"20",x"49",x"2F",x"4F",x"20",x"6F", -- 0x3FB8
		x"6E",x"6C",x"79",x"00",x"46",x"69",x"6C",x"65", -- 0x3FC0
		x"20",x"6E",x"6F",x"74",x"20",x"4F",x"50",x"45", -- 0x3FC8
		x"4E",x"00",x"20",x"69",x"6E",x"20",x"00",x"4F", -- 0x3FD0
		x"6B",x"0D",x"0A",x"00",x"42",x"72",x"65",x"61", -- 0x3FD8
		x"6B",x"00",x"21",x"04",x"00",x"39",x"7E",x"23", -- 0x3FE0
		x"FE",x"82",x"C0",x"4E",x"23",x"46",x"23",x"E5", -- 0x3FE8
		x"60",x"69",x"7A",x"B3",x"EB",x"28",x"02",x"EB", -- 0x3FF0
		x"E7",x"01",x"16",x"00",x"E1",x"C8",x"09",x"18", -- 0x3FF8
		x"E5",x"CD",x"39",x"54",x"44",x"4D",x"ED",x"78", -- 0x4000
		x"C3",x"CF",x"4F",x"CD",x"2F",x"54",x"D5",x"CF", -- 0x4008
		x"2C",x"CD",x"1C",x"52",x"C1",x"C9",x"CD",x"0B", -- 0x4010
		x"40",x"ED",x"79",x"C9",x"CD",x"0B",x"40",x"C5", -- 0x4018
		x"F5",x"1E",x"00",x"2B",x"D7",x"28",x"05",x"CF", -- 0x4020
		x"2C",x"CD",x"1C",x"52",x"F1",x"57",x"C1",x"CD", -- 0x4028
		x"BD",x"00",x"ED",x"78",x"AB",x"A2",x"28",x"F7", -- 0x4030
		x"C9",x"CD",x"F8",x"FE",x"2A",x"1C",x"F4",x"7C", -- 0x4038
		x"A5",x"3C",x"28",x"08",x"3A",x"BB",x"F6",x"B7", -- 0x4040
		x"1E",x"15",x"20",x"23",x"C3",x"01",x"64",x"2A", -- 0x4048
		x"A3",x"F6",x"22",x"1C",x"F4",x"1E",x"02",x"01", -- 0x4050
		x"1E",x"0B",x"01",x"1E",x"01",x"01",x"1E",x"0A", -- 0x4058
		x"01",x"1E",x"12",x"01",x"1E",x"16",x"01",x"1E", -- 0x4060
		x"06",x"01",x"1E",x"18",x"01",x"1E",x"0D",x"CD", -- 0x4068
		x"B1",x"FF",x"AF",x"32",x"7C",x"F8",x"2A",x"19", -- 0x4070
		x"F4",x"7C",x"B5",x"28",x"0A",x"3A",x"1B",x"F4", -- 0x4078
		x"77",x"21",x"00",x"00",x"22",x"19",x"F4",x"FB", -- 0x4080
		x"2A",x"1C",x"F4",x"22",x"B3",x"F6",x"7C",x"A5", -- 0x4088
		x"3C",x"28",x"03",x"22",x"B5",x"F6",x"01",x"A4", -- 0x4090
		x"40",x"18",x"03",x"01",x"1E",x"41",x"2A",x"B1", -- 0x4098
		x"F6",x"C3",x"F0",x"62",x"C1",x"7B",x"4B",x"32", -- 0x40A0
		x"14",x"F4",x"2A",x"AF",x"F6",x"22",x"B7",x"F6", -- 0x40A8
		x"EB",x"2A",x"B3",x"F6",x"7C",x"A5",x"3C",x"28", -- 0x40B0
		x"07",x"22",x"BE",x"F6",x"EB",x"22",x"C0",x"F6", -- 0x40B8
		x"2A",x"B9",x"F6",x"7C",x"B5",x"EB",x"21",x"BB", -- 0x40C0
		x"F6",x"28",x"08",x"A6",x"20",x"05",x"35",x"EB", -- 0x40C8
		x"C3",x"20",x"46",x"AF",x"77",x"59",x"CD",x"23", -- 0x40D0
		x"73",x"21",x"75",x"3D",x"CD",x"FD",x"FE",x"7B", -- 0x40D8
		x"FE",x"3C",x"30",x"08",x"FE",x"32",x"30",x"06", -- 0x40E0
		x"FE",x"1A",x"38",x"05",x"3E",x"2F",x"D6",x"18", -- 0x40E8
		x"5F",x"CD",x"5D",x"48",x"23",x"1D",x"20",x"F9", -- 0x40F0
		x"E5",x"2A",x"B3",x"F6",x"E3",x"CD",x"02",x"FF", -- 0x40F8
		x"E5",x"CD",x"D2",x"00",x"E1",x"7E",x"FE",x"3F", -- 0x4100
		x"20",x"06",x"E1",x"21",x"75",x"3D",x"18",x"DC", -- 0x4108
		x"3E",x"07",x"DF",x"CD",x"78",x"66",x"E1",x"7C", -- 0x4110
		x"A5",x"3C",x"C4",x"0A",x"34",x"3E",x"C1",x"CD", -- 0x4118
		x"D2",x"00",x"CD",x"04",x"73",x"CD",x"7B",x"6D", -- 0x4120
		x"CD",x"07",x"FF",x"CD",x"23",x"73",x"21",x"D7", -- 0x4128
		x"3F",x"CD",x"78",x"66",x"CD",x"0C",x"FF",x"21", -- 0x4130
		x"FF",x"FF",x"22",x"1C",x"F4",x"21",x"0F",x"F4", -- 0x4138
		x"22",x"AF",x"F6",x"3A",x"AA",x"F6",x"B7",x"28", -- 0x4140
		x"16",x"2A",x"AB",x"F6",x"E5",x"CD",x"12",x"34", -- 0x4148
		x"D1",x"D5",x"CD",x"95",x"42",x"3E",x"2A",x"38", -- 0x4150
		x"02",x"3E",x"20",x"DF",x"32",x"AA",x"F6",x"CD", -- 0x4158
		x"4A",x"01",x"20",x"0C",x"CD",x"AE",x"00",x"30", -- 0x4160
		x"0A",x"AF",x"32",x"AA",x"F6",x"C3",x"34",x"41", -- 0x4168
		x"CD",x"74",x"73",x"D7",x"3C",x"3D",x"28",x"BC", -- 0x4170
		x"F5",x"CD",x"69",x"47",x"30",x"06",x"CD",x"4A", -- 0x4178
		x"01",x"CA",x"55",x"40",x"CD",x"14",x"45",x"3A", -- 0x4180
		x"AA",x"F6",x"B7",x"28",x"08",x"FE",x"2A",x"20", -- 0x4188
		x"04",x"BE",x"20",x"01",x"23",x"7A",x"B3",x"28", -- 0x4190
		x"06",x"7E",x"FE",x"20",x"20",x"01",x"23",x"D5", -- 0x4198
		x"CD",x"B2",x"42",x"D1",x"F1",x"22",x"AF",x"F6", -- 0x41A0
		x"CD",x"11",x"FF",x"38",x"07",x"AF",x"32",x"AA", -- 0x41A8
		x"F6",x"C3",x"48",x"6D",x"D5",x"C5",x"D7",x"B7", -- 0x41B0
		x"F5",x"3A",x"AA",x"F6",x"A7",x"28",x"03",x"F1", -- 0x41B8
		x"37",x"F5",x"ED",x"53",x"B5",x"F6",x"2A",x"AD", -- 0x41C0
		x"F6",x"19",x"38",x"0B",x"D5",x"11",x"FA",x"FF", -- 0x41C8
		x"E7",x"D1",x"22",x"AB",x"F6",x"38",x"04",x"AF", -- 0x41D0
		x"32",x"AA",x"F6",x"CD",x"95",x"42",x"38",x"0D", -- 0x41D8
		x"F1",x"F5",x"20",x"06",x"D2",x"1C",x"48",x"C5", -- 0x41E0
		x"18",x"4D",x"B7",x"18",x"07",x"F1",x"F5",x"20", -- 0x41E8
		x"02",x"38",x"F4",x"37",x"C5",x"F5",x"E5",x"CD", -- 0x41F0
		x"EA",x"54",x"E1",x"F1",x"C1",x"C5",x"DC",x"05", -- 0x41F8
		x"54",x"D1",x"F1",x"D5",x"28",x"31",x"D1",x"21", -- 0x4200
		x"00",x"00",x"22",x"B9",x"F6",x"2A",x"C2",x"F6", -- 0x4208
		x"E3",x"C1",x"E5",x"09",x"E5",x"CD",x"50",x"62", -- 0x4210
		x"E1",x"22",x"C2",x"F6",x"EB",x"74",x"C1",x"D1", -- 0x4218
		x"E5",x"23",x"23",x"73",x"23",x"72",x"23",x"11", -- 0x4220
		x"1F",x"F4",x"0B",x"0B",x"0B",x"0B",x"1A",x"77", -- 0x4228
		x"23",x"13",x"0B",x"79",x"B0",x"20",x"F7",x"CD", -- 0x4230
		x"16",x"FF",x"D1",x"CD",x"57",x"42",x"2A",x"64", -- 0x4238
		x"F8",x"22",x"BC",x"F6",x"CD",x"9A",x"62",x"CD", -- 0x4240
		x"1B",x"FF",x"2A",x"BC",x"F6",x"22",x"64",x"F8", -- 0x4248
		x"C3",x"34",x"41",x"2A",x"76",x"F6",x"EB",x"62", -- 0x4250
		x"6B",x"7E",x"23",x"B6",x"C8",x"23",x"23",x"23", -- 0x4258
		x"7E",x"B7",x"28",x"0E",x"FE",x"20",x"30",x"F7", -- 0x4260
		x"FE",x"0B",x"38",x"F3",x"CD",x"6A",x"46",x"D7", -- 0x4268
		x"18",x"EF",x"23",x"EB",x"73",x"23",x"72",x"18", -- 0x4270
		x"DE",x"11",x"00",x"00",x"D5",x"28",x"09",x"D1", -- 0x4278
		x"CD",x"5F",x"47",x"D5",x"28",x"0B",x"CF",x"F2", -- 0x4280
		x"11",x"FA",x"FF",x"C4",x"5F",x"47",x"C2",x"55", -- 0x4288
		x"40",x"EB",x"D1",x"E3",x"E5",x"2A",x"76",x"F6", -- 0x4290
		x"44",x"4D",x"7E",x"23",x"B6",x"2B",x"C8",x"23", -- 0x4298
		x"23",x"7E",x"23",x"66",x"6F",x"E7",x"60",x"69", -- 0x42A0
		x"7E",x"23",x"66",x"6F",x"3F",x"C8",x"3F",x"D0", -- 0x42A8
		x"18",x"E6",x"AF",x"32",x"65",x"F6",x"32",x"64", -- 0x42B0
		x"F6",x"CD",x"20",x"FF",x"01",x"3B",x"01",x"11", -- 0x42B8
		x"1F",x"F4",x"7E",x"B7",x"20",x"13",x"21",x"40", -- 0x42C0
		x"01",x"7D",x"91",x"4F",x"7C",x"98",x"47",x"21", -- 0x42C8
		x"1E",x"F4",x"AF",x"12",x"13",x"12",x"13",x"12", -- 0x42D0
		x"C9",x"FE",x"22",x"CA",x"16",x"43",x"FE",x"20", -- 0x42D8
		x"28",x"07",x"3A",x"64",x"F6",x"B7",x"7E",x"28", -- 0x42E0
		x"3D",x"23",x"F5",x"FE",x"01",x"20",x"04",x"7E", -- 0x42E8
		x"A7",x"3E",x"01",x"C4",x"E0",x"44",x"F1",x"D6", -- 0x42F0
		x"3A",x"28",x"06",x"FE",x"4A",x"20",x"08",x"3E", -- 0x42F8
		x"01",x"32",x"64",x"F6",x"32",x"65",x"F6",x"D6", -- 0x4300
		x"55",x"20",x"B7",x"F5",x"7E",x"B7",x"E3",x"7C", -- 0x4308
		x"E1",x"28",x"B3",x"BE",x"28",x"D3",x"F5",x"7E", -- 0x4310
		x"23",x"FE",x"01",x"20",x"04",x"7E",x"A7",x"3E", -- 0x4318
		x"01",x"C4",x"E0",x"44",x"18",x"E6",x"23",x"B7", -- 0x4320
		x"FA",x"C2",x"42",x"FE",x"01",x"20",x"07",x"7E", -- 0x4328
		x"A7",x"28",x"93",x"23",x"18",x"8C",x"2B",x"FE", -- 0x4330
		x"3F",x"3E",x"91",x"D5",x"C5",x"CA",x"A3",x"43", -- 0x4338
		x"7E",x"FE",x"5F",x"CA",x"A3",x"43",x"11",x"26", -- 0x4340
		x"3D",x"CD",x"A9",x"4E",x"CD",x"A8",x"64",x"DA", -- 0x4348
		x"1D",x"44",x"E5",x"CD",x"25",x"FF",x"21",x"3E", -- 0x4350
		x"3A",x"D6",x"41",x"87",x"4F",x"06",x"00",x"09", -- 0x4358
		x"5E",x"23",x"56",x"E1",x"23",x"E5",x"CD",x"A9", -- 0x4360
		x"4E",x"4F",x"1A",x"E6",x"7F",x"CA",x"EB",x"44", -- 0x4368
		x"23",x"B9",x"20",x"24",x"1A",x"13",x"B7",x"F2", -- 0x4370
		x"66",x"43",x"F1",x"1A",x"CD",x"2A",x"FF",x"B7", -- 0x4378
		x"FA",x"A2",x"43",x"C1",x"D1",x"F6",x"80",x"F5", -- 0x4380
		x"3E",x"FF",x"CD",x"E0",x"44",x"AF",x"32",x"65", -- 0x4388
		x"F6",x"F1",x"CD",x"E0",x"44",x"C3",x"C2",x"42", -- 0x4390
		x"E1",x"1A",x"13",x"B7",x"F2",x"99",x"43",x"13", -- 0x4398
		x"18",x"C3",x"2B",x"F5",x"CD",x"2F",x"FF",x"11", -- 0x43A0
		x"B5",x"43",x"4F",x"1A",x"B7",x"28",x"15",x"13", -- 0x43A8
		x"B9",x"20",x"F8",x"18",x"11",x"8C",x"A9",x"AA", -- 0x43B0
		x"A8",x"A7",x"E1",x"A1",x"8A",x"93",x"9E",x"89", -- 0x43B8
		x"8E",x"DA",x"8D",x"00",x"AF",x"C2",x"3E",x"01", -- 0x43C0
		x"32",x"65",x"F6",x"F1",x"C1",x"D1",x"FE",x"A1", -- 0x43C8
		x"F5",x"CC",x"DE",x"44",x"F1",x"FE",x"CA",x"28", -- 0x43D0
		x"04",x"FE",x"5F",x"20",x"29",x"D4",x"E0",x"44", -- 0x43D8
		x"23",x"CD",x"A9",x"4E",x"A7",x"CA",x"C6",x"42", -- 0x43E0
		x"FA",x"E0",x"43",x"FE",x"01",x"20",x"07",x"23", -- 0x43E8
		x"7E",x"A7",x"28",x"F1",x"18",x"EA",x"FE",x"20", -- 0x43F0
		x"28",x"E3",x"FE",x"3A",x"28",x"3C",x"FE",x"28", -- 0x43F8
		x"28",x"38",x"FE",x"30",x"18",x"D7",x"FE",x"E6", -- 0x4400
		x"C2",x"B4",x"44",x"F5",x"CD",x"DE",x"44",x"3E", -- 0x4408
		x"8F",x"CD",x"E0",x"44",x"F1",x"E5",x"21",x"00", -- 0x4410
		x"00",x"E3",x"C3",x"18",x"43",x"7E",x"FE",x"2E", -- 0x4418
		x"28",x"0A",x"FE",x"3A",x"D2",x"A2",x"44",x"FE", -- 0x4420
		x"30",x"DA",x"A2",x"44",x"3A",x"65",x"F6",x"B7", -- 0x4428
		x"7E",x"C1",x"D1",x"FA",x"E9",x"42",x"28",x"1F", -- 0x4430
		x"FE",x"2E",x"CA",x"E9",x"42",x"3E",x"0E",x"CD", -- 0x4438
		x"E0",x"44",x"D5",x"CD",x"69",x"47",x"CD",x"14", -- 0x4440
		x"45",x"E3",x"EB",x"7D",x"CD",x"E0",x"44",x"7C", -- 0x4448
		x"E1",x"CD",x"E0",x"44",x"C3",x"C2",x"42",x"D5", -- 0x4450
		x"C5",x"7E",x"CD",x"99",x"32",x"CD",x"14",x"45", -- 0x4458
		x"C1",x"D1",x"E5",x"3A",x"63",x"F6",x"FE",x"02", -- 0x4460
		x"20",x"15",x"2A",x"F8",x"F7",x"7C",x"B7",x"3E", -- 0x4468
		x"02",x"20",x"0C",x"7D",x"65",x"2E",x"0F",x"FE", -- 0x4470
		x"0A",x"30",x"D0",x"C6",x"11",x"18",x"D1",x"F5", -- 0x4478
		x"0F",x"C6",x"1B",x"CD",x"E0",x"44",x"21",x"F6", -- 0x4480
		x"F7",x"3A",x"63",x"F6",x"FE",x"02",x"20",x"03", -- 0x4488
		x"21",x"F8",x"F7",x"F1",x"F5",x"7E",x"CD",x"E0", -- 0x4490
		x"44",x"F1",x"23",x"3D",x"20",x"F6",x"E1",x"C3", -- 0x4498
		x"C2",x"42",x"11",x"25",x"3D",x"13",x"1A",x"E6", -- 0x44A0
		x"7F",x"CA",x"FA",x"44",x"13",x"BE",x"1A",x"20", -- 0x44A8
		x"F4",x"C3",x"09",x"45",x"FE",x"26",x"C2",x"E9", -- 0x44B0
		x"42",x"E5",x"D7",x"E1",x"CD",x"AA",x"4E",x"FE", -- 0x44B8
		x"48",x"28",x"0D",x"FE",x"4F",x"28",x"05",x"3E", -- 0x44C0
		x"26",x"C3",x"E9",x"42",x"3E",x"0B",x"18",x"02", -- 0x44C8
		x"3E",x"0C",x"CD",x"E0",x"44",x"D5",x"C5",x"CD", -- 0x44D0
		x"B8",x"4E",x"C1",x"C3",x"49",x"44",x"3E",x"3A", -- 0x44D8
		x"12",x"13",x"0B",x"79",x"B0",x"C0",x"1E",x"19", -- 0x44E0
		x"C3",x"6F",x"40",x"CD",x"34",x"FF",x"E1",x"2B", -- 0x44E8
		x"3D",x"32",x"65",x"F6",x"CD",x"A9",x"4E",x"C3", -- 0x44F0
		x"CC",x"43",x"7E",x"FE",x"20",x"30",x"0A",x"FE", -- 0x44F8
		x"09",x"28",x"06",x"FE",x"0A",x"28",x"02",x"3E", -- 0x4500
		x"20",x"F5",x"3A",x"65",x"F6",x"3C",x"28",x"01", -- 0x4508
		x"3D",x"C3",x"C8",x"43",x"2B",x"7E",x"FE",x"20", -- 0x4510
		x"28",x"FA",x"FE",x"09",x"28",x"F6",x"FE",x"0A", -- 0x4518
		x"28",x"F2",x"23",x"C9",x"3E",x"64",x"32",x"A5", -- 0x4520
		x"F6",x"CD",x"80",x"48",x"C1",x"E5",x"CD",x"5B", -- 0x4528
		x"48",x"22",x"A1",x"F6",x"21",x"02",x"00",x"39", -- 0x4530
		x"CD",x"E6",x"3F",x"20",x"17",x"09",x"D5",x"2B", -- 0x4538
		x"56",x"2B",x"5E",x"23",x"23",x"E5",x"2A",x"A1", -- 0x4540
		x"F6",x"E7",x"E1",x"D1",x"20",x"EA",x"D1",x"F9", -- 0x4548
		x"22",x"B1",x"F6",x"0E",x"D1",x"EB",x"0E",x"0C", -- 0x4550
		x"CD",x"5E",x"62",x"E5",x"2A",x"A1",x"F6",x"E3", -- 0x4558
		x"E5",x"2A",x"1C",x"F4",x"E3",x"CF",x"D9",x"EF", -- 0x4560
		x"CA",x"6D",x"40",x"F5",x"CD",x"64",x"4C",x"F1", -- 0x4568
		x"E5",x"30",x"18",x"F2",x"C2",x"45",x"CD",x"8A", -- 0x4570
		x"2F",x"E3",x"11",x"01",x"00",x"7E",x"FE",x"DC", -- 0x4578
		x"CC",x"0E",x"52",x"D5",x"E5",x"EB",x"CD",x"AB", -- 0x4580
		x"2E",x"18",x"5D",x"CD",x"3A",x"30",x"D1",x"21", -- 0x4588
		x"F8",x"FF",x"39",x"F9",x"D5",x"CD",x"10",x"2F", -- 0x4590
		x"E1",x"7E",x"FE",x"DC",x"11",x"1B",x"2D",x"3E", -- 0x4598
		x"01",x"20",x"0F",x"D7",x"CD",x"64",x"4C",x"E5", -- 0x45A0
		x"CD",x"3A",x"30",x"CD",x"71",x"2E",x"11",x"F6", -- 0x45A8
		x"F7",x"E1",x"44",x"4D",x"21",x"F8",x"FF",x"39", -- 0x45B0
		x"F9",x"F5",x"C5",x"CD",x"F3",x"2E",x"E1",x"F1", -- 0x45B8
		x"18",x"2D",x"CD",x"B2",x"2F",x"CD",x"CC",x"2E", -- 0x45C0
		x"E1",x"C5",x"D5",x"01",x"41",x"10",x"11",x"00", -- 0x45C8
		x"00",x"CD",x"39",x"FF",x"7E",x"FE",x"DC",x"3E", -- 0x45D0
		x"01",x"20",x"0E",x"CD",x"65",x"4C",x"E5",x"CD", -- 0x45D8
		x"B2",x"2F",x"CD",x"CC",x"2E",x"CD",x"71",x"2E", -- 0x45E0
		x"E1",x"D5",x"C5",x"C5",x"C5",x"C5",x"C5",x"B7", -- 0x45E8
		x"20",x"02",x"3E",x"02",x"4F",x"EF",x"47",x"C5", -- 0x45F0
		x"E5",x"2A",x"A7",x"F6",x"E3",x"06",x"82",x"C5", -- 0x45F8
		x"33",x"CD",x"3E",x"FF",x"ED",x"73",x"B1",x"F6", -- 0x4600
		x"CD",x"BA",x"00",x"3A",x"D8",x"FB",x"B7",x"C4", -- 0x4608
		x"89",x"63",x"FB",x"22",x"AF",x"F6",x"7E",x"FE", -- 0x4610
		x"3A",x"28",x"25",x"B7",x"C2",x"55",x"40",x"23", -- 0x4618
		x"7E",x"23",x"B6",x"CA",x"39",x"40",x"23",x"5E", -- 0x4620
		x"23",x"56",x"EB",x"22",x"1C",x"F4",x"3A",x"C4", -- 0x4628
		x"F7",x"B7",x"28",x"0B",x"D5",x"3E",x"5B",x"DF", -- 0x4630
		x"CD",x"12",x"34",x"3E",x"5D",x"DF",x"D1",x"EB", -- 0x4638
		x"D7",x"11",x"01",x"46",x"D5",x"C8",x"CD",x"43", -- 0x4640
		x"FF",x"FE",x"5F",x"CA",x"A7",x"55",x"D6",x"81", -- 0x4648
		x"DA",x"80",x"48",x"FE",x"58",x"D2",x"AD",x"51", -- 0x4650
		x"07",x"4F",x"06",x"00",x"EB",x"21",x"2E",x"39", -- 0x4658
		x"09",x"4E",x"23",x"46",x"C5",x"EB",x"CD",x"48", -- 0x4660
		x"FF",x"23",x"7E",x"FE",x"3A",x"D0",x"FE",x"20", -- 0x4668
		x"28",x"F4",x"30",x"6C",x"B7",x"C8",x"FE",x"0B", -- 0x4670
		x"38",x"61",x"FE",x"1E",x"20",x"05",x"3A",x"68", -- 0x4678
		x"F6",x"B7",x"C9",x"FE",x"10",x"28",x"34",x"F5", -- 0x4680
		x"23",x"32",x"68",x"F6",x"D6",x"1C",x"30",x"30", -- 0x4688
		x"D6",x"F5",x"30",x"06",x"FE",x"FE",x"20",x"16", -- 0x4690
		x"7E",x"23",x"22",x"66",x"F6",x"26",x"00",x"6F", -- 0x4698
		x"22",x"6A",x"F6",x"3E",x"02",x"32",x"69",x"F6", -- 0x46A0
		x"21",x"E6",x"46",x"F1",x"B7",x"C9",x"7E",x"23", -- 0x46A8
		x"23",x"22",x"66",x"F6",x"2B",x"66",x"18",x"E7", -- 0x46B0
		x"CD",x"E8",x"46",x"2A",x"66",x"F6",x"18",x"AA", -- 0x46B8
		x"3C",x"07",x"32",x"69",x"F6",x"D5",x"C5",x"11", -- 0x46C0
		x"6A",x"F6",x"EB",x"47",x"CD",x"F7",x"2E",x"EB", -- 0x46C8
		x"C1",x"D1",x"22",x"66",x"F6",x"F1",x"21",x"E6", -- 0x46D0
		x"46",x"B7",x"C9",x"FE",x"09",x"D2",x"66",x"46", -- 0x46D8
		x"FE",x"30",x"3F",x"3C",x"3D",x"C9",x"1E",x"10", -- 0x46E0
		x"3A",x"68",x"F6",x"FE",x"0F",x"30",x"13",x"FE", -- 0x46E8
		x"0D",x"38",x"0F",x"2A",x"6A",x"F6",x"20",x"07", -- 0x46F0
		x"23",x"23",x"23",x"5E",x"23",x"56",x"EB",x"C3", -- 0x46F8
		x"36",x"32",x"3A",x"69",x"F6",x"32",x"63",x"F6", -- 0x4700
		x"FE",x"02",x"20",x"06",x"2A",x"6A",x"F6",x"22", -- 0x4708
		x"F8",x"F7",x"21",x"6A",x"F6",x"C3",x"08",x"2F", -- 0x4710
		x"1E",x"03",x"01",x"1E",x"02",x"01",x"1E",x"04", -- 0x4718
		x"01",x"1E",x"08",x"CD",x"A7",x"64",x"01",x"55", -- 0x4720
		x"40",x"C5",x"D8",x"D6",x"41",x"4F",x"47",x"D7", -- 0x4728
		x"FE",x"F2",x"20",x"09",x"D7",x"CD",x"A7",x"64", -- 0x4730
		x"D8",x"D6",x"41",x"47",x"D7",x"78",x"91",x"D8", -- 0x4738
		x"3C",x"E3",x"21",x"CA",x"F6",x"06",x"00",x"09", -- 0x4740
		x"73",x"23",x"3D",x"20",x"FB",x"E1",x"7E",x"FE", -- 0x4748
		x"2C",x"C0",x"D7",x"18",x"CE",x"D7",x"CD",x"0F", -- 0x4750
		x"52",x"F0",x"1E",x"05",x"C3",x"6F",x"40",x"7E", -- 0x4758
		x"FE",x"2E",x"ED",x"5B",x"B5",x"F6",x"CA",x"66", -- 0x4760
		x"46",x"2B",x"D7",x"FE",x"0E",x"28",x"02",x"FE", -- 0x4768
		x"0D",x"ED",x"5B",x"6A",x"F6",x"CA",x"66",x"46", -- 0x4770
		x"AF",x"32",x"68",x"F6",x"11",x"00",x"00",x"2B", -- 0x4778
		x"D7",x"D0",x"E5",x"F5",x"21",x"98",x"19",x"E7", -- 0x4780
		x"38",x"11",x"62",x"6B",x"19",x"29",x"19",x"29", -- 0x4788
		x"F1",x"D6",x"30",x"5F",x"16",x"00",x"19",x"EB", -- 0x4790
		x"E1",x"18",x"E5",x"F1",x"E1",x"C9",x"CA",x"9A", -- 0x4798
		x"62",x"FE",x"0E",x"28",x"05",x"FE",x"0D",x"C2", -- 0x47A0
		x"5B",x"6B",x"CD",x"A1",x"62",x"01",x"01",x"46", -- 0x47A8
		x"18",x"35",x"0E",x"03",x"CD",x"5E",x"62",x"CD", -- 0x47B0
		x"69",x"47",x"C1",x"E5",x"E5",x"2A",x"1C",x"F4", -- 0x47B8
		x"E3",x"01",x"00",x"00",x"C5",x"01",x"01",x"46", -- 0x47C0
		x"3E",x"8D",x"F5",x"33",x"C5",x"18",x"1C",x"E5", -- 0x47C8
		x"E5",x"2A",x"1C",x"F4",x"E3",x"C5",x"3E",x"8D", -- 0x47D0
		x"F5",x"33",x"EB",x"2B",x"22",x"AF",x"F6",x"23", -- 0x47D8
		x"ED",x"73",x"B1",x"F6",x"C3",x"20",x"46",x"C5", -- 0x47E0
		x"CD",x"69",x"47",x"3A",x"68",x"F6",x"FE",x"0D", -- 0x47E8
		x"EB",x"C8",x"FE",x"0E",x"C2",x"55",x"40",x"EB", -- 0x47F0
		x"E5",x"2A",x"66",x"F6",x"E3",x"CD",x"5D",x"48", -- 0x47F8
		x"23",x"E5",x"2A",x"1C",x"F4",x"E7",x"E1",x"DC", -- 0x4800
		x"98",x"42",x"D4",x"95",x"42",x"30",x"0D",x"0B", -- 0x4808
		x"3E",x"0D",x"32",x"A9",x"F6",x"E1",x"CD",x"83", -- 0x4810
		x"55",x"60",x"69",x"C9",x"1E",x"08",x"C3",x"6F", -- 0x4818
		x"40",x"CD",x"4D",x"FF",x"22",x"A7",x"F6",x"16", -- 0x4820
		x"FF",x"CD",x"E2",x"3F",x"FE",x"8D",x"28",x"01", -- 0x4828
		x"2B",x"F9",x"22",x"B1",x"F6",x"1E",x"03",x"C2", -- 0x4830
		x"6F",x"40",x"E1",x"7C",x"B5",x"28",x"06",x"7E", -- 0x4838
		x"E6",x"01",x"C4",x"3E",x"63",x"C1",x"21",x"01", -- 0x4840
		x"46",x"E3",x"EB",x"2A",x"A7",x"F6",x"2B",x"D7", -- 0x4848
		x"C2",x"E8",x"47",x"60",x"69",x"22",x"1C",x"F4", -- 0x4850
		x"EB",x"3E",x"E1",x"01",x"3A",x"0E",x"00",x"06", -- 0x4858
		x"00",x"79",x"48",x"47",x"2B",x"D7",x"B7",x"C8", -- 0x4860
		x"B8",x"C8",x"23",x"FE",x"22",x"28",x"F2",x"3C", -- 0x4868
		x"28",x"F3",x"D6",x"8C",x"20",x"EE",x"B8",x"8A", -- 0x4870
		x"57",x"18",x"E9",x"F1",x"C6",x"03",x"18",x"12", -- 0x4878
		x"CD",x"A4",x"5E",x"CF",x"EF",x"ED",x"53",x"A7", -- 0x4880
		x"F6",x"D5",x"3A",x"63",x"F6",x"F5",x"CD",x"64", -- 0x4888
		x"4C",x"F1",x"E3",x"47",x"3A",x"63",x"F6",x"B8", -- 0x4890
		x"78",x"28",x"06",x"CD",x"7A",x"51",x"3A",x"63", -- 0x4898
		x"F6",x"11",x"F6",x"F7",x"FE",x"02",x"20",x"03", -- 0x48A0
		x"11",x"F8",x"F7",x"E5",x"FE",x"03",x"20",x"2E", -- 0x48A8
		x"2A",x"F8",x"F7",x"E5",x"23",x"5E",x"23",x"56", -- 0x48B0
		x"21",x"1E",x"F4",x"E7",x"38",x"14",x"2A",x"C6", -- 0x48B8
		x"F6",x"E7",x"D1",x"30",x"15",x"21",x"97",x"F6", -- 0x48C0
		x"E7",x"38",x"06",x"21",x"79",x"F6",x"E7",x"38", -- 0x48C8
		x"09",x"3E",x"D1",x"CD",x"EE",x"67",x"EB",x"CD", -- 0x48D0
		x"11",x"66",x"CD",x"EE",x"67",x"E3",x"CD",x"F3", -- 0x48D8
		x"2E",x"D1",x"E1",x"C9",x"FE",x"A6",x"20",x"25", -- 0x48E0
		x"D7",x"CF",x"89",x"CD",x"69",x"47",x"7A",x"B3", -- 0x48E8
		x"28",x"09",x"CD",x"93",x"42",x"50",x"59",x"E1", -- 0x48F0
		x"D2",x"1C",x"48",x"ED",x"53",x"B9",x"F6",x"D8", -- 0x48F8
		x"3A",x"BB",x"F6",x"B7",x"7B",x"C8",x"3A",x"14", -- 0x4900
		x"F4",x"5F",x"C3",x"96",x"40",x"CD",x"10",x"78", -- 0x4908
		x"38",x"31",x"C5",x"D7",x"CF",x"8D",x"AF",x"C1", -- 0x4910
		x"C5",x"B9",x"D2",x"55",x"40",x"F5",x"CD",x"69", -- 0x4918
		x"47",x"7A",x"B3",x"28",x"09",x"CD",x"93",x"42", -- 0x4920
		x"50",x"59",x"E1",x"D2",x"1C",x"48",x"F1",x"C1", -- 0x4928
		x"F5",x"80",x"C5",x"CD",x"5C",x"78",x"2B",x"D7", -- 0x4930
		x"C1",x"D1",x"C8",x"C5",x"D5",x"CF",x"2C",x"F1", -- 0x4938
		x"3C",x"18",x"D4",x"CD",x"1C",x"52",x"7E",x"47", -- 0x4940
		x"FE",x"8D",x"28",x"03",x"CF",x"89",x"2B",x"4B", -- 0x4948
		x"0D",x"78",x"CA",x"46",x"46",x"CD",x"6A",x"47", -- 0x4950
		x"FE",x"2C",x"C0",x"18",x"F3",x"3A",x"BB",x"F6", -- 0x4958
		x"B7",x"20",x"09",x"32",x"B9",x"F6",x"32",x"BA", -- 0x4960
		x"F6",x"C3",x"64",x"40",x"3C",x"32",x"14",x"F4", -- 0x4968
		x"7E",x"FE",x"83",x"28",x"10",x"CD",x"69",x"47", -- 0x4970
		x"C0",x"7A",x"B3",x"28",x"0C",x"CD",x"EB",x"47", -- 0x4978
		x"AF",x"32",x"BB",x"F6",x"C9",x"D7",x"C0",x"18", -- 0x4980
		x"05",x"AF",x"32",x"BB",x"F6",x"3C",x"2A",x"B7", -- 0x4988
		x"F6",x"EB",x"2A",x"B3",x"F6",x"22",x"1C",x"F4", -- 0x4990
		x"EB",x"C0",x"7E",x"B7",x"20",x"04",x"23",x"23", -- 0x4998
		x"23",x"23",x"23",x"AF",x"32",x"BB",x"F6",x"C3", -- 0x49A0
		x"5B",x"48",x"CD",x"1C",x"52",x"C0",x"B7",x"CA", -- 0x49A8
		x"5A",x"47",x"C3",x"6F",x"40",x"11",x"0A",x"00", -- 0x49B0
		x"D5",x"28",x"16",x"CD",x"5F",x"47",x"EB",x"E3", -- 0x49B8
		x"28",x"10",x"EB",x"CF",x"2C",x"ED",x"5B",x"AD", -- 0x49C0
		x"F6",x"28",x"06",x"CD",x"69",x"47",x"C2",x"55", -- 0x49C8
		x"40",x"EB",x"7C",x"B5",x"CA",x"5A",x"47",x"22", -- 0x49D0
		x"AD",x"F6",x"32",x"AA",x"F6",x"E1",x"22",x"AB", -- 0x49D8
		x"F6",x"C1",x"C3",x"34",x"41",x"CD",x"64",x"4C", -- 0x49E0
		x"7E",x"FE",x"2C",x"CC",x"66",x"46",x"FE",x"89", -- 0x49E8
		x"28",x"03",x"CF",x"DA",x"2B",x"E5",x"CD",x"A1", -- 0x49F0
		x"2E",x"E1",x"28",x"10",x"D7",x"C8",x"FE",x"0E", -- 0x49F8
		x"CA",x"E8",x"47",x"FE",x"0D",x"C2",x"46",x"46", -- 0x4A00
		x"2A",x"6A",x"F6",x"C9",x"16",x"01",x"CD",x"5B", -- 0x4A08
		x"48",x"B7",x"C8",x"D7",x"FE",x"A1",x"20",x"F6", -- 0x4A10
		x"15",x"20",x"F3",x"18",x"DF",x"3E",x"01",x"32", -- 0x4A18
		x"16",x"F4",x"18",x"05",x"0E",x"02",x"CD",x"57", -- 0x4A20
		x"6D",x"2B",x"D7",x"CC",x"28",x"73",x"CA",x"FF", -- 0x4A28
		x"4A",x"FE",x"E4",x"CA",x"B1",x"60",x"FE",x"DB", -- 0x4A30
		x"CA",x"C6",x"4A",x"FE",x"DF",x"CA",x"C6",x"4A", -- 0x4A38
		x"E5",x"FE",x"2C",x"28",x"4F",x"FE",x"3B",x"CA", -- 0x4A40
		x"FA",x"4A",x"C1",x"CD",x"64",x"4C",x"E5",x"EF", -- 0x4A48
		x"28",x"3B",x"CD",x"25",x"34",x"CD",x"35",x"66", -- 0x4A50
		x"36",x"20",x"2A",x"F8",x"F7",x"34",x"CD",x"52", -- 0x4A58
		x"FF",x"CD",x"4A",x"01",x"20",x"23",x"2A",x"F8", -- 0x4A60
		x"F7",x"3A",x"16",x"F4",x"B7",x"28",x"08",x"3A", -- 0x4A68
		x"15",x"F4",x"86",x"FE",x"FF",x"18",x"0A",x"3A", -- 0x4A70
		x"B0",x"F3",x"47",x"3A",x"61",x"F6",x"86",x"3D", -- 0x4A78
		x"B8",x"38",x"06",x"CC",x"31",x"73",x"C4",x"28", -- 0x4A80
		x"73",x"CD",x"7B",x"66",x"B7",x"CC",x"7B",x"66", -- 0x4A88
		x"E1",x"C3",x"29",x"4A",x"CD",x"57",x"FF",x"01", -- 0x4A90
		x"08",x"00",x"2A",x"64",x"F8",x"09",x"CD",x"4A", -- 0x4A98
		x"01",x"7E",x"20",x"1B",x"3A",x"16",x"F4",x"B7", -- 0x4AA0
		x"28",x"07",x"3A",x"15",x"F4",x"FE",x"EE",x"18", -- 0x4AA8
		x"08",x"3A",x"B2",x"F3",x"47",x"3A",x"61",x"F6", -- 0x4AB0
		x"B8",x"D4",x"28",x"73",x"D2",x"FA",x"4A",x"D6", -- 0x4AB8
		x"0E",x"30",x"FC",x"2F",x"18",x"2D",x"F5",x"CD", -- 0x4AC0
		x"1B",x"52",x"CF",x"29",x"2B",x"F1",x"D6",x"DF", -- 0x4AC8
		x"E5",x"28",x"1C",x"01",x"08",x"00",x"2A",x"64", -- 0x4AD0
		x"F8",x"09",x"CD",x"4A",x"01",x"7E",x"20",x"0F", -- 0x4AD8
		x"3A",x"16",x"F4",x"B7",x"CA",x"EC",x"4A",x"3A", -- 0x4AE0
		x"15",x"F4",x"18",x"03",x"3A",x"61",x"F6",x"2F", -- 0x4AE8
		x"83",x"30",x"07",x"3C",x"47",x"3E",x"20",x"DF", -- 0x4AF0
		x"10",x"FD",x"E1",x"D7",x"C3",x"2E",x"4A",x"CD", -- 0x4AF8
		x"5C",x"FF",x"AF",x"32",x"16",x"F4",x"E5",x"67", -- 0x4B00
		x"6F",x"22",x"64",x"F8",x"E1",x"C9",x"FE",x"85", -- 0x4B08
		x"C2",x"A7",x"58",x"CF",x"85",x"FE",x"23",x"CA", -- 0x4B10
		x"8F",x"6D",x"CD",x"7B",x"4B",x"CD",x"A4",x"5E", -- 0x4B18
		x"CD",x"58",x"30",x"D5",x"E5",x"CD",x"B1",x"00", -- 0x4B20
		x"D1",x"C1",x"DA",x"FE",x"63",x"C5",x"D5",x"06", -- 0x4B28
		x"00",x"CD",x"38",x"66",x"E1",x"3E",x"03",x"C3", -- 0x4B30
		x"92",x"48",x"3F",x"52",x"65",x"64",x"6F",x"20", -- 0x4B38
		x"66",x"72",x"6F",x"6D",x"20",x"73",x"74",x"61", -- 0x4B40
		x"72",x"74",x"0D",x"0A",x"00",x"CD",x"61",x"FF", -- 0x4B48
		x"3A",x"A6",x"F6",x"B7",x"C2",x"4F",x"40",x"C1", -- 0x4B50
		x"21",x"3A",x"4B",x"CD",x"78",x"66",x"2A",x"AF", -- 0x4B58
		x"F6",x"C9",x"CD",x"55",x"6D",x"E5",x"21",x"5D", -- 0x4B60
		x"F5",x"C3",x"9B",x"4B",x"FE",x"23",x"28",x"F2", -- 0x4B68
		x"E5",x"F5",x"CD",x"D2",x"00",x"F1",x"E1",x"01", -- 0x4B70
		x"8B",x"4B",x"C5",x"FE",x"22",x"3E",x"00",x"C0", -- 0x4B78
		x"CD",x"36",x"66",x"CF",x"3B",x"E5",x"CD",x"7B", -- 0x4B80
		x"66",x"E1",x"C9",x"E5",x"CD",x"B4",x"00",x"C1", -- 0x4B88
		x"DA",x"FE",x"63",x"23",x"7E",x"B7",x"2B",x"C5", -- 0x4B90
		x"CA",x"5A",x"48",x"36",x"2C",x"18",x"05",x"E5", -- 0x4B98
		x"2A",x"C8",x"F6",x"F6",x"AF",x"32",x"A6",x"F6", -- 0x4BA0
		x"E3",x"01",x"CF",x"2C",x"CD",x"A4",x"5E",x"E3", -- 0x4BA8
		x"D5",x"7E",x"FE",x"2C",x"28",x"1B",x"3A",x"A6", -- 0x4BB0
		x"F6",x"B7",x"C2",x"40",x"4C",x"3E",x"3F",x"DF", -- 0x4BB8
		x"CD",x"B4",x"00",x"D1",x"C1",x"DA",x"FE",x"63", -- 0x4BC0
		x"23",x"7E",x"2B",x"B7",x"C5",x"CA",x"5A",x"48", -- 0x4BC8
		x"D5",x"CD",x"4A",x"01",x"C2",x"83",x"6D",x"EF", -- 0x4BD0
		x"F5",x"20",x"22",x"D7",x"57",x"47",x"FE",x"22", -- 0x4BD8
		x"28",x"0C",x"3A",x"A6",x"F6",x"B7",x"57",x"28", -- 0x4BE0
		x"02",x"16",x"3A",x"06",x"2C",x"2B",x"CD",x"39", -- 0x4BE8
		x"66",x"F1",x"C6",x"03",x"EB",x"21",x"05",x"4C", -- 0x4BF0
		x"E3",x"D5",x"C3",x"93",x"48",x"D7",x"01",x"F1", -- 0x4BF8
		x"4B",x"C5",x"C3",x"99",x"32",x"2B",x"D7",x"28", -- 0x4C00
		x"05",x"FE",x"2C",x"C2",x"4D",x"4B",x"E3",x"2B", -- 0x4C08
		x"D7",x"C2",x"AA",x"4B",x"D1",x"3A",x"A6",x"F6", -- 0x4C10
		x"B7",x"EB",x"C2",x"DE",x"63",x"D5",x"CD",x"4A", -- 0x4C18
		x"01",x"20",x"08",x"7E",x"B7",x"21",x"2F",x"4C", -- 0x4C20
		x"C4",x"78",x"66",x"E1",x"C3",x"FF",x"4A",x"3F", -- 0x4C28
		x"45",x"78",x"74",x"72",x"61",x"20",x"69",x"67", -- 0x4C30
		x"6E",x"6F",x"72",x"65",x"64",x"0D",x"0A",x"00", -- 0x4C38
		x"CD",x"5B",x"48",x"B7",x"20",x"11",x"23",x"7E", -- 0x4C40
		x"23",x"B6",x"1E",x"04",x"CA",x"6F",x"40",x"23", -- 0x4C48
		x"5E",x"23",x"56",x"ED",x"53",x"A3",x"F6",x"D7", -- 0x4C50
		x"FE",x"84",x"20",x"E4",x"C3",x"D1",x"4B",x"CF", -- 0x4C58
		x"EF",x"01",x"CF",x"28",x"2B",x"16",x"00",x"D5", -- 0x4C60
		x"0E",x"01",x"CD",x"5E",x"62",x"CD",x"66",x"FF", -- 0x4C68
		x"CD",x"C7",x"4D",x"22",x"BC",x"F6",x"2A",x"BC", -- 0x4C70
		x"F6",x"C1",x"7E",x"22",x"9D",x"F6",x"FE",x"EE", -- 0x4C78
		x"D8",x"FE",x"F1",x"38",x"5F",x"D6",x"F1",x"5F", -- 0x4C80
		x"20",x"09",x"3A",x"63",x"F6",x"FE",x"03",x"7B", -- 0x4C88
		x"CA",x"87",x"67",x"FE",x"0C",x"D0",x"21",x"3B", -- 0x4C90
		x"3D",x"16",x"00",x"19",x"78",x"56",x"BA",x"D0", -- 0x4C98
		x"C5",x"01",x"76",x"4C",x"C5",x"7A",x"CD",x"6B", -- 0x4CA0
		x"FF",x"FE",x"51",x"38",x"50",x"E6",x"FE",x"FE", -- 0x4CA8
		x"7A",x"28",x"4A",x"21",x"F8",x"F7",x"3A",x"63", -- 0x4CB0
		x"F6",x"D6",x"03",x"CA",x"6D",x"40",x"B7",x"2A", -- 0x4CB8
		x"F8",x"F7",x"E5",x"FA",x"D5",x"4C",x"2A",x"F6", -- 0x4CC0
		x"F7",x"E5",x"E2",x"D5",x"4C",x"2A",x"FC",x"F7", -- 0x4CC8
		x"E5",x"2A",x"FA",x"F7",x"E5",x"C6",x"03",x"4B", -- 0x4CD0
		x"47",x"C5",x"01",x"22",x"4D",x"C5",x"2A",x"9D", -- 0x4CD8
		x"F6",x"C3",x"67",x"4C",x"16",x"00",x"D6",x"EE", -- 0x4CE0
		x"38",x"1E",x"FE",x"03",x"30",x"1A",x"FE",x"01", -- 0x4CE8
		x"17",x"AA",x"BA",x"57",x"DA",x"55",x"40",x"22", -- 0x4CF0
		x"9D",x"F6",x"D7",x"18",x"E9",x"D5",x"CD",x"8A", -- 0x4CF8
		x"2F",x"D1",x"E5",x"01",x"78",x"4F",x"18",x"D5", -- 0x4D00
		x"78",x"FE",x"64",x"D0",x"C5",x"D5",x"11",x"05", -- 0x4D08
		x"64",x"21",x"57",x"4F",x"E5",x"EF",x"C2",x"B3", -- 0x4D10
		x"4C",x"2A",x"F8",x"F7",x"E5",x"01",x"C8",x"65", -- 0x4D18
		x"18",x"BB",x"C1",x"79",x"32",x"64",x"F6",x"3A", -- 0x4D20
		x"63",x"F6",x"B8",x"20",x"0B",x"FE",x"02",x"28", -- 0x4D28
		x"1F",x"FE",x"04",x"CA",x"9D",x"4D",x"30",x"2B", -- 0x4D30
		x"57",x"78",x"FE",x"08",x"28",x"22",x"7A",x"FE", -- 0x4D38
		x"08",x"28",x"44",x"78",x"FE",x"04",x"28",x"52", -- 0x4D40
		x"7A",x"FE",x"03",x"CA",x"6D",x"40",x"30",x"54", -- 0x4D48
		x"21",x"69",x"3D",x"06",x"00",x"09",x"09",x"4E", -- 0x4D50
		x"23",x"46",x"D1",x"2A",x"F8",x"F7",x"C5",x"C9", -- 0x4D58
		x"CD",x"3A",x"30",x"CD",x"0D",x"2F",x"E1",x"22", -- 0x4D60
		x"FA",x"F7",x"E1",x"22",x"FC",x"F7",x"C1",x"D1", -- 0x4D68
		x"CD",x"C1",x"2E",x"CD",x"3A",x"30",x"21",x"51", -- 0x4D70
		x"3D",x"3A",x"64",x"F6",x"07",x"85",x"6F",x"8C", -- 0x4D78
		x"95",x"67",x"7E",x"23",x"66",x"6F",x"E9",x"78", -- 0x4D80
		x"F5",x"CD",x"0D",x"2F",x"F1",x"32",x"63",x"F6", -- 0x4D88
		x"FE",x"04",x"28",x"DA",x"E1",x"22",x"F8",x"F7", -- 0x4D90
		x"18",x"D9",x"CD",x"B2",x"2F",x"C1",x"D1",x"21", -- 0x4D98
		x"5D",x"3D",x"18",x"D5",x"E1",x"CD",x"B1",x"2E", -- 0x4DA0
		x"CD",x"CB",x"2F",x"CD",x"CC",x"2E",x"E1",x"22", -- 0x4DA8
		x"F6",x"F7",x"E1",x"22",x"F8",x"F7",x"18",x"E7", -- 0x4DB0
		x"E5",x"EB",x"CD",x"CB",x"2F",x"E1",x"CD",x"B1", -- 0x4DB8
		x"2E",x"CD",x"CB",x"2F",x"C3",x"65",x"32",x"D7", -- 0x4DC0
		x"CA",x"6A",x"40",x"DA",x"99",x"32",x"CD",x"A8", -- 0x4DC8
		x"64",x"D2",x"9B",x"4E",x"FE",x"20",x"DA",x"B8", -- 0x4DD0
		x"46",x"CD",x"70",x"FF",x"3C",x"CA",x"FC",x"4E", -- 0x4DD8
		x"3D",x"FE",x"F1",x"28",x"E2",x"FE",x"F2",x"CA", -- 0x4DE0
		x"8D",x"4E",x"FE",x"22",x"CA",x"36",x"66",x"FE", -- 0x4DE8
		x"E0",x"CA",x"63",x"4F",x"FE",x"26",x"CA",x"B8", -- 0x4DF0
		x"4E",x"FE",x"E2",x"20",x"0A",x"D7",x"3A",x"14", -- 0x4DF8
		x"F4",x"E5",x"CD",x"CF",x"4F",x"E1",x"C9",x"FE", -- 0x4E00
		x"E1",x"20",x"0A",x"D7",x"E5",x"2A",x"B3",x"F6", -- 0x4E08
		x"CD",x"36",x"32",x"E1",x"C9",x"FE",x"ED",x"CA", -- 0x4E10
		x"03",x"58",x"FE",x"CB",x"CA",x"00",x"79",x"FE", -- 0x4E18
		x"C7",x"CA",x"84",x"7A",x"FE",x"C8",x"CA",x"47", -- 0x4E20
		x"7B",x"FE",x"C9",x"CA",x"CB",x"7B",x"FE",x"C1", -- 0x4E28
		x"CA",x"1B",x"79",x"FE",x"EA",x"CA",x"3E",x"7C", -- 0x4E30
		x"FE",x"E9",x"CA",x"43",x"7C",x"FE",x"E7",x"20", -- 0x4E38
		x"23",x"D7",x"CF",x"28",x"FE",x"23",x"20",x"0B", -- 0x4E40
		x"CD",x"1B",x"52",x"E5",x"CD",x"6D",x"6A",x"EB", -- 0x4E48
		x"E1",x"18",x"03",x"CD",x"5D",x"5F",x"CF",x"29", -- 0x4E50
		x"E5",x"EB",x"7C",x"B5",x"CA",x"5A",x"47",x"CD", -- 0x4E58
		x"99",x"2F",x"E1",x"C9",x"FE",x"DD",x"CA",x"D5", -- 0x4E60
		x"4F",x"FE",x"E5",x"CA",x"EB",x"68",x"FE",x"EC", -- 0x4E68
		x"CA",x"47",x"73",x"FE",x"E3",x"CA",x"29",x"68", -- 0x4E70
		x"FE",x"85",x"CA",x"87",x"6C",x"FE",x"E8",x"CA", -- 0x4E78
		x"0A",x"79",x"FE",x"DE",x"CA",x"40",x"50",x"CD", -- 0x4E80
		x"62",x"4C",x"CF",x"29",x"C9",x"16",x"7D",x"CD", -- 0x4E88
		x"67",x"4C",x"2A",x"BC",x"F6",x"E5",x"CD",x"86", -- 0x4E90
		x"2E",x"E1",x"C9",x"CD",x"A4",x"5E",x"E5",x"EB", -- 0x4E98
		x"22",x"F8",x"F7",x"EF",x"C4",x"08",x"2F",x"E1", -- 0x4EA0
		x"C9",x"7E",x"FE",x"61",x"D8",x"FE",x"7B",x"D0", -- 0x4EA8
		x"E6",x"5F",x"C9",x"FE",x"26",x"C2",x"69",x"47", -- 0x4EB0
		x"11",x"00",x"00",x"D7",x"CD",x"AA",x"4E",x"01", -- 0x4EB8
		x"02",x"01",x"FE",x"42",x"28",x"0F",x"01",x"08", -- 0x4EC0
		x"03",x"FE",x"4F",x"28",x"08",x"01",x"10",x"04", -- 0x4EC8
		x"FE",x"48",x"C2",x"55",x"40",x"23",x"7E",x"EB", -- 0x4ED0
		x"CD",x"AA",x"4E",x"FE",x"3A",x"38",x"06",x"FE", -- 0x4ED8
		x"41",x"38",x"14",x"D6",x"07",x"D6",x"30",x"B9", -- 0x4EE0
		x"30",x"0D",x"C5",x"29",x"DA",x"67",x"40",x"10", -- 0x4EE8
		x"FA",x"C1",x"B5",x"6F",x"EB",x"18",x"DE",x"CD", -- 0x4EF0
		x"99",x"2F",x"EB",x"C9",x"23",x"7E",x"D6",x"81", -- 0x4EF8
		x"06",x"00",x"07",x"4F",x"C5",x"D7",x"79",x"FE", -- 0x4F00
		x"05",x"30",x"16",x"CD",x"62",x"4C",x"CF",x"2C", -- 0x4F08
		x"CD",x"58",x"30",x"EB",x"2A",x"F8",x"F7",x"E3", -- 0x4F10
		x"E5",x"EB",x"CD",x"1C",x"52",x"EB",x"E3",x"18", -- 0x4F18
		x"1A",x"CD",x"87",x"4E",x"E3",x"7D",x"FE",x"0C", -- 0x4F20
		x"38",x"0D",x"FE",x"1B",x"CD",x"75",x"FF",x"30", -- 0x4F28
		x"06",x"EF",x"E5",x"DC",x"3A",x"30",x"E1",x"11", -- 0x4F30
		x"99",x"4E",x"D5",x"01",x"DE",x"39",x"CD",x"7A", -- 0x4F38
		x"FF",x"09",x"4E",x"23",x"66",x"69",x"E9",x"15", -- 0x4F40
		x"FE",x"F2",x"C8",x"FE",x"2D",x"C8",x"14",x"FE", -- 0x4F48
		x"2B",x"C8",x"FE",x"F1",x"C8",x"2B",x"C9",x"3C", -- 0x4F50
		x"8F",x"C1",x"A0",x"C6",x"FF",x"9F",x"CD",x"9A", -- 0x4F58
		x"2E",x"18",x"12",x"16",x"5A",x"CD",x"67",x"4C", -- 0x4F60
		x"CD",x"8A",x"2F",x"7D",x"2F",x"6F",x"7C",x"2F", -- 0x4F68
		x"67",x"22",x"F8",x"F7",x"C1",x"C3",x"76",x"4C", -- 0x4F70
		x"78",x"F5",x"CD",x"8A",x"2F",x"F1",x"D1",x"FE", -- 0x4F78
		x"7A",x"CA",x"3A",x"32",x"FE",x"7B",x"CA",x"E6", -- 0x4F80
		x"31",x"01",x"D1",x"4F",x"C5",x"FE",x"46",x"20", -- 0x4F88
		x"06",x"7B",x"B5",x"6F",x"7C",x"B2",x"C9",x"FE", -- 0x4F90
		x"50",x"20",x"06",x"7B",x"A5",x"6F",x"7C",x"A2", -- 0x4F98
		x"C9",x"FE",x"3C",x"20",x"06",x"7B",x"AD",x"6F", -- 0x4FA0
		x"7C",x"AA",x"C9",x"FE",x"32",x"20",x"08",x"7B", -- 0x4FA8
		x"AD",x"2F",x"6F",x"7C",x"AA",x"2F",x"C9",x"7D", -- 0x4FB0
		x"2F",x"A3",x"2F",x"6F",x"7C",x"2F",x"A2",x"2F", -- 0x4FB8
		x"C9",x"B7",x"ED",x"52",x"C3",x"36",x"32",x"3A", -- 0x4FC0
		x"15",x"F4",x"18",x"03",x"3A",x"61",x"F6",x"6F", -- 0x4FC8
		x"AF",x"67",x"C3",x"99",x"2F",x"CD",x"F4",x"4F", -- 0x4FD0
		x"D5",x"CD",x"87",x"4E",x"E3",x"5E",x"23",x"56", -- 0x4FD8
		x"21",x"97",x"32",x"E5",x"D5",x"3A",x"63",x"F6", -- 0x4FE0
		x"F5",x"FE",x"03",x"CC",x"D3",x"67",x"F1",x"EB", -- 0x4FE8
		x"21",x"F6",x"F7",x"C9",x"D7",x"01",x"00",x"00", -- 0x4FF0
		x"FE",x"1B",x"30",x"0B",x"FE",x"11",x"38",x"07", -- 0x4FF8
		x"D7",x"3A",x"6A",x"F6",x"B7",x"17",x"4F",x"EB", -- 0x5000
		x"21",x"9A",x"F3",x"09",x"EB",x"C9",x"CD",x"F4", -- 0x5008
		x"4F",x"D5",x"CF",x"EF",x"CD",x"2F",x"54",x"E3", -- 0x5010
		x"73",x"23",x"72",x"E1",x"C9",x"FE",x"DD",x"28", -- 0x5018
		x"ED",x"CD",x"A1",x"51",x"CD",x"93",x"51",x"EB", -- 0x5020
		x"73",x"23",x"72",x"EB",x"7E",x"FE",x"28",x"C2", -- 0x5028
		x"5B",x"48",x"D7",x"CD",x"A4",x"5E",x"7E",x"FE", -- 0x5030
		x"29",x"CA",x"5B",x"48",x"CF",x"2C",x"18",x"F3", -- 0x5038
		x"CD",x"A1",x"51",x"3A",x"63",x"F6",x"B7",x"F5", -- 0x5040
		x"22",x"BC",x"F6",x"EB",x"7E",x"23",x"66",x"6F", -- 0x5048
		x"7C",x"B5",x"CA",x"61",x"40",x"7E",x"FE",x"28", -- 0x5050
		x"C2",x"F4",x"50",x"D7",x"22",x"9D",x"F6",x"EB", -- 0x5058
		x"2A",x"BC",x"F6",x"CF",x"28",x"AF",x"F5",x"E5", -- 0x5060
		x"EB",x"3E",x"80",x"32",x"A5",x"F6",x"CD",x"A4", -- 0x5068
		x"5E",x"EB",x"E3",x"3A",x"63",x"F6",x"F5",x"D5", -- 0x5070
		x"CD",x"64",x"4C",x"22",x"BC",x"F6",x"E1",x"22", -- 0x5078
		x"9D",x"F6",x"F1",x"CD",x"7A",x"51",x"0E",x"04", -- 0x5080
		x"CD",x"5E",x"62",x"21",x"F8",x"FF",x"39",x"F9", -- 0x5088
		x"CD",x"10",x"2F",x"3A",x"63",x"F6",x"F5",x"2A", -- 0x5090
		x"BC",x"F6",x"7E",x"FE",x"29",x"28",x"0E",x"CF", -- 0x5098
		x"2C",x"E5",x"2A",x"9D",x"F6",x"CF",x"2C",x"18", -- 0x50A0
		x"C0",x"F1",x"32",x"4E",x"F7",x"F1",x"B7",x"28", -- 0x50A8
		x"38",x"32",x"63",x"F6",x"21",x"00",x"00",x"39", -- 0x50B0
		x"CD",x"08",x"2F",x"21",x"08",x"00",x"39",x"F9", -- 0x50B8
		x"D1",x"2E",x"03",x"1B",x"1B",x"1B",x"3A",x"63", -- 0x50C0
		x"F6",x"85",x"47",x"3A",x"4E",x"F7",x"4F",x"80", -- 0x50C8
		x"FE",x"64",x"D2",x"5A",x"47",x"F5",x"7D",x"06", -- 0x50D0
		x"00",x"21",x"50",x"F7",x"09",x"4F",x"CD",x"8E", -- 0x50D8
		x"51",x"01",x"A9",x"50",x"C5",x"C5",x"C3",x"9E", -- 0x50E0
		x"48",x"2A",x"BC",x"F6",x"D7",x"E5",x"2A",x"9D", -- 0x50E8
		x"F6",x"CF",x"29",x"3E",x"D5",x"22",x"9D",x"F6", -- 0x50F0
		x"3A",x"E6",x"F6",x"C6",x"04",x"F5",x"0F",x"4F", -- 0x50F8
		x"CD",x"5E",x"62",x"F1",x"4F",x"2F",x"3C",x"6F", -- 0x5100
		x"26",x"FF",x"39",x"F9",x"E5",x"11",x"E4",x"F6", -- 0x5108
		x"CD",x"8E",x"51",x"E1",x"22",x"E4",x"F6",x"2A", -- 0x5110
		x"4E",x"F7",x"22",x"E6",x"F6",x"44",x"4D",x"21", -- 0x5118
		x"E8",x"F6",x"11",x"50",x"F7",x"CD",x"8E",x"51", -- 0x5120
		x"67",x"6F",x"22",x"4E",x"F7",x"2A",x"BA",x"F7", -- 0x5128
		x"23",x"22",x"BA",x"F7",x"7C",x"B5",x"32",x"B7", -- 0x5130
		x"F7",x"2A",x"9D",x"F6",x"CD",x"5F",x"4C",x"2B", -- 0x5138
		x"D7",x"C2",x"55",x"40",x"EF",x"20",x"0F",x"11", -- 0x5140
		x"98",x"F6",x"2A",x"F8",x"F7",x"E7",x"38",x"06", -- 0x5148
		x"CD",x"11",x"66",x"CD",x"58",x"66",x"2A",x"E4", -- 0x5150
		x"F6",x"54",x"5D",x"23",x"23",x"4E",x"23",x"46", -- 0x5158
		x"03",x"03",x"03",x"03",x"21",x"E4",x"F6",x"CD", -- 0x5160
		x"8E",x"51",x"EB",x"F9",x"2A",x"BA",x"F7",x"2B", -- 0x5168
		x"22",x"BA",x"F7",x"7C",x"B5",x"32",x"B7",x"F7", -- 0x5170
		x"E1",x"F1",x"E5",x"E6",x"07",x"21",x"47",x"3D", -- 0x5178
		x"4F",x"06",x"00",x"09",x"CD",x"41",x"4F",x"E1", -- 0x5180
		x"C9",x"1A",x"77",x"23",x"13",x"0B",x"78",x"B1", -- 0x5188
		x"20",x"F7",x"C9",x"E5",x"2A",x"1C",x"F4",x"23", -- 0x5190
		x"7C",x"B5",x"E1",x"C0",x"1E",x"0C",x"C3",x"6F", -- 0x5198
		x"40",x"CF",x"DE",x"3E",x"80",x"32",x"A5",x"F6", -- 0x51A0
		x"B6",x"4F",x"C3",x"A9",x"5E",x"FE",x"7E",x"20", -- 0x51A8
		x"15",x"23",x"7E",x"23",x"FE",x"83",x"CA",x"6E", -- 0x51B0
		x"69",x"FE",x"A3",x"CA",x"BF",x"77",x"FE",x"85", -- 0x51B8
		x"CA",x"B1",x"77",x"CD",x"7F",x"FF",x"C3",x"55", -- 0x51C0
		x"40",x"CD",x"1C",x"52",x"CD",x"84",x"FF",x"A7", -- 0x51C8
		x"28",x"0D",x"3A",x"B0",x"FC",x"A7",x"7B",x"28", -- 0x51D0
		x"04",x"FE",x"21",x"30",x"02",x"FE",x"29",x"D2", -- 0x51D8
		x"5A",x"47",x"3A",x"B0",x"F3",x"BB",x"C8",x"3E", -- 0x51E0
		x"0C",x"DF",x"7B",x"32",x"B0",x"F3",x"3A",x"B0", -- 0x51E8
		x"FC",x"3D",x"7B",x"20",x"05",x"32",x"AF",x"F3", -- 0x51F0
		x"18",x"03",x"32",x"AE",x"F3",x"3E",x"0C",x"DF", -- 0x51F8
		x"7B",x"D6",x"0E",x"30",x"FC",x"C6",x"1C",x"2F", -- 0x5200
		x"3C",x"83",x"32",x"B2",x"F3",x"C9",x"D7",x"CD", -- 0x5208
		x"64",x"4C",x"E5",x"CD",x"8A",x"2F",x"EB",x"E1", -- 0x5210
		x"7A",x"B7",x"C9",x"D7",x"CD",x"64",x"4C",x"CD", -- 0x5218
		x"12",x"52",x"C2",x"5A",x"47",x"2B",x"D7",x"7B", -- 0x5220
		x"C9",x"3E",x"01",x"32",x"16",x"F4",x"CD",x"89", -- 0x5228
		x"FF",x"C1",x"CD",x"79",x"42",x"C5",x"21",x"FF", -- 0x5230
		x"FF",x"22",x"1C",x"F4",x"E1",x"D1",x"4E",x"23", -- 0x5238
		x"46",x"23",x"78",x"B1",x"CA",x"1F",x"41",x"CD", -- 0x5240
		x"4A",x"01",x"CC",x"BA",x"00",x"C5",x"4E",x"23", -- 0x5248
		x"46",x"23",x"C5",x"E3",x"EB",x"E7",x"C1",x"DA", -- 0x5250
		x"1E",x"41",x"E3",x"E5",x"C5",x"EB",x"22",x"B5", -- 0x5258
		x"F6",x"CD",x"12",x"34",x"E1",x"7E",x"FE",x"09", -- 0x5260
		x"28",x"03",x"3E",x"20",x"DF",x"CD",x"84",x"52", -- 0x5268
		x"21",x"5E",x"F5",x"CD",x"7B",x"52",x"CD",x"28", -- 0x5270
		x"73",x"18",x"BB",x"7E",x"B7",x"C8",x"CD",x"67", -- 0x5278
		x"73",x"23",x"18",x"F7",x"01",x"5E",x"F5",x"16", -- 0x5280
		x"FF",x"AF",x"32",x"64",x"F6",x"18",x"04",x"03", -- 0x5288
		x"23",x"15",x"C8",x"7E",x"B7",x"02",x"C8",x"FE", -- 0x5290
		x"0B",x"38",x"25",x"FE",x"20",x"DA",x"61",x"53", -- 0x5298
		x"FE",x"22",x"20",x"0A",x"3A",x"64",x"F6",x"EE", -- 0x52A0
		x"01",x"32",x"64",x"F6",x"3E",x"22",x"FE",x"3A", -- 0x52A8
		x"20",x"0E",x"3A",x"64",x"F6",x"1F",x"38",x"06", -- 0x52B0
		x"17",x"E6",x"FD",x"32",x"64",x"F6",x"3E",x"3A", -- 0x52B8
		x"B7",x"F2",x"8F",x"52",x"3A",x"64",x"F6",x"1F", -- 0x52C0
		x"38",x"2E",x"1F",x"1F",x"30",x"3E",x"7E",x"FE", -- 0x52C8
		x"E6",x"E5",x"C5",x"21",x"F5",x"52",x"E5",x"C0", -- 0x52D0
		x"0B",x"0A",x"FE",x"4D",x"C0",x"0B",x"0A",x"FE", -- 0x52D8
		x"45",x"C0",x"0B",x"0A",x"FE",x"52",x"C0",x"0B", -- 0x52E0
		x"0A",x"FE",x"3A",x"C0",x"F1",x"F1",x"E1",x"14", -- 0x52E8
		x"14",x"14",x"14",x"18",x"25",x"C1",x"E1",x"7E", -- 0x52F0
		x"C3",x"8F",x"52",x"3A",x"64",x"F6",x"F6",x"02", -- 0x52F8
		x"32",x"64",x"F6",x"AF",x"C9",x"3A",x"64",x"F6", -- 0x5300
		x"F6",x"04",x"18",x"F4",x"17",x"38",x"E9",x"7E", -- 0x5308
		x"FE",x"84",x"CC",x"FB",x"52",x"FE",x"8F",x"CC", -- 0x5310
		x"05",x"53",x"7E",x"3C",x"7E",x"20",x"04",x"23", -- 0x5318
		x"7E",x"E6",x"7F",x"23",x"FE",x"A1",x"20",x"02", -- 0x5320
		x"0B",x"14",x"E5",x"C5",x"D5",x"CD",x"8E",x"FF", -- 0x5328
		x"21",x"71",x"3A",x"47",x"0E",x"40",x"0C",x"23", -- 0x5330
		x"54",x"5D",x"7E",x"B7",x"28",x"F8",x"23",x"F2", -- 0x5338
		x"3A",x"53",x"7E",x"B8",x"20",x"F1",x"EB",x"79", -- 0x5340
		x"D1",x"C1",x"FE",x"5B",x"20",x"02",x"7E",x"23", -- 0x5348
		x"5F",x"E6",x"7F",x"02",x"03",x"15",x"CA",x"A7", -- 0x5350
		x"66",x"B3",x"F2",x"4E",x"53",x"E1",x"C3",x"93", -- 0x5358
		x"52",x"2B",x"D7",x"D5",x"C5",x"F5",x"CD",x"E8", -- 0x5360
		x"46",x"F1",x"01",x"7E",x"53",x"C5",x"FE",x"0B", -- 0x5368
		x"CA",x"1E",x"37",x"FE",x"0C",x"CA",x"22",x"37", -- 0x5370
		x"2A",x"6A",x"F6",x"C3",x"25",x"34",x"C1",x"D1", -- 0x5378
		x"3A",x"68",x"F6",x"1E",x"4F",x"FE",x"0B",x"28", -- 0x5380
		x"06",x"FE",x"0C",x"1E",x"48",x"20",x"0B",x"3E", -- 0x5388
		x"26",x"02",x"03",x"15",x"C8",x"7B",x"02",x"03", -- 0x5390
		x"15",x"C8",x"3A",x"69",x"F6",x"FE",x"04",x"1E", -- 0x5398
		x"00",x"38",x"06",x"1E",x"21",x"28",x"02",x"1E", -- 0x53A0
		x"23",x"7E",x"FE",x"20",x"20",x"01",x"23",x"7E", -- 0x53A8
		x"23",x"B7",x"28",x"20",x"02",x"03",x"15",x"C8", -- 0x53B0
		x"3A",x"69",x"F6",x"FE",x"04",x"38",x"F0",x"0B", -- 0x53B8
		x"0A",x"03",x"20",x"04",x"FE",x"2E",x"28",x"08", -- 0x53C0
		x"FE",x"44",x"28",x"04",x"FE",x"45",x"20",x"DF", -- 0x53C8
		x"1E",x"00",x"18",x"DB",x"7B",x"B7",x"28",x"04", -- 0x53D0
		x"02",x"03",x"15",x"C8",x"2A",x"66",x"F6",x"C3", -- 0x53D8
		x"93",x"52",x"CD",x"79",x"42",x"C5",x"CD",x"EA", -- 0x53E0
		x"54",x"C1",x"D1",x"C5",x"C5",x"CD",x"95",x"42", -- 0x53E8
		x"30",x"05",x"54",x"5D",x"E3",x"E5",x"E7",x"D2", -- 0x53F0
		x"5A",x"47",x"21",x"D7",x"3F",x"CD",x"78",x"66", -- 0x53F8
		x"C1",x"21",x"37",x"42",x"E3",x"EB",x"2A",x"C2", -- 0x5400
		x"F6",x"1A",x"02",x"03",x"13",x"E7",x"20",x"F9", -- 0x5408
		x"60",x"69",x"22",x"C2",x"F6",x"22",x"C4",x"F6", -- 0x5410
		x"22",x"C6",x"F6",x"C9",x"CD",x"39",x"54",x"7E", -- 0x5418
		x"C3",x"CF",x"4F",x"CD",x"2F",x"54",x"D5",x"CF", -- 0x5420
		x"2C",x"CD",x"1C",x"52",x"D1",x"12",x"C9",x"CD", -- 0x5428
		x"64",x"4C",x"E5",x"CD",x"39",x"54",x"EB",x"E1", -- 0x5430
		x"C9",x"01",x"8A",x"2F",x"C5",x"EF",x"F8",x"CD", -- 0x5438
		x"93",x"FF",x"CD",x"71",x"2E",x"F8",x"CD",x"B2", -- 0x5440
		x"2F",x"01",x"45",x"32",x"11",x"76",x"80",x"CD", -- 0x5448
		x"21",x"2F",x"D8",x"01",x"45",x"65",x"11",x"53", -- 0x5450
		x"60",x"CD",x"21",x"2F",x"D2",x"67",x"40",x"01", -- 0x5458
		x"C5",x"65",x"11",x"53",x"60",x"C3",x"4E",x"32", -- 0x5460
		x"01",x"0A",x"00",x"C5",x"50",x"58",x"28",x"26", -- 0x5468
		x"FE",x"2C",x"28",x"09",x"D5",x"CD",x"5F",x"47", -- 0x5470
		x"42",x"4B",x"D1",x"28",x"19",x"CF",x"2C",x"CD", -- 0x5478
		x"5F",x"47",x"28",x"12",x"F1",x"CF",x"2C",x"D5", -- 0x5480
		x"CD",x"69",x"47",x"C2",x"55",x"40",x"7A",x"B3", -- 0x5488
		x"CA",x"5A",x"47",x"EB",x"E3",x"EB",x"C5",x"CD", -- 0x5490
		x"95",x"42",x"D1",x"D5",x"C5",x"CD",x"95",x"42", -- 0x5498
		x"60",x"69",x"D1",x"E7",x"EB",x"DA",x"5A",x"47", -- 0x54A0
		x"D1",x"C1",x"F1",x"E5",x"D5",x"18",x"0E",x"09", -- 0x54A8
		x"DA",x"5A",x"47",x"EB",x"E5",x"21",x"F9",x"FF", -- 0x54B0
		x"E7",x"E1",x"DA",x"5A",x"47",x"D5",x"5E",x"23", -- 0x54B8
		x"56",x"7A",x"B3",x"EB",x"D1",x"28",x"07",x"7E", -- 0x54C0
		x"23",x"B6",x"2B",x"EB",x"20",x"E1",x"C5",x"CD", -- 0x54C8
		x"F6",x"54",x"C1",x"D1",x"E1",x"D5",x"5E",x"23", -- 0x54D0
		x"56",x"7A",x"B3",x"28",x"14",x"EB",x"E3",x"EB", -- 0x54D8
		x"23",x"73",x"23",x"72",x"EB",x"09",x"EB",x"E1", -- 0x54E0
		x"18",x"EB",x"3A",x"A9",x"F6",x"B7",x"C8",x"18", -- 0x54E8
		x"06",x"01",x"1E",x"41",x"C5",x"FE",x"F6",x"AF", -- 0x54F0
		x"32",x"A9",x"F6",x"2A",x"76",x"F6",x"2B",x"23", -- 0x54F8
		x"7E",x"23",x"B6",x"C8",x"23",x"5E",x"23",x"56", -- 0x5500
		x"D7",x"B7",x"28",x"F3",x"4F",x"3A",x"A9",x"F6", -- 0x5508
		x"B7",x"79",x"28",x"56",x"CD",x"98",x"FF",x"FE", -- 0x5510
		x"A6",x"20",x"14",x"D7",x"FE",x"89",x"20",x"E9", -- 0x5518
		x"D7",x"FE",x"0E",x"20",x"E4",x"D5",x"CD",x"71", -- 0x5520
		x"47",x"7A",x"B3",x"20",x"0A",x"18",x"27",x"FE", -- 0x5528
		x"0E",x"20",x"D5",x"D5",x"CD",x"71",x"47",x"E5", -- 0x5530
		x"CD",x"95",x"42",x"0B",x"3E",x"0D",x"38",x"3C", -- 0x5538
		x"CD",x"23",x"73",x"21",x"5A",x"55",x"D5",x"CD", -- 0x5540
		x"78",x"66",x"E1",x"CD",x"12",x"34",x"C1",x"E1", -- 0x5548
		x"E5",x"C5",x"CD",x"0A",x"34",x"E1",x"D1",x"2B", -- 0x5550
		x"18",x"AE",x"55",x"6E",x"64",x"65",x"66",x"69", -- 0x5558
		x"6E",x"65",x"64",x"20",x"6C",x"69",x"6E",x"65", -- 0x5560
		x"20",x"00",x"FE",x"0D",x"20",x"EA",x"D5",x"CD", -- 0x5568
		x"71",x"47",x"E5",x"EB",x"23",x"23",x"23",x"4E", -- 0x5570
		x"23",x"46",x"3E",x"0E",x"21",x"55",x"55",x"E5", -- 0x5578
		x"2A",x"66",x"F6",x"E5",x"2B",x"70",x"2B",x"71", -- 0x5580
		x"2B",x"77",x"E1",x"C9",x"7E",x"E3",x"BE",x"23", -- 0x5588
		x"E3",x"C2",x"55",x"40",x"C3",x"66",x"46",x"3A", -- 0x5590
		x"63",x"F6",x"FE",x"08",x"30",x"05",x"D6",x"03", -- 0x5598
		x"B7",x"37",x"C9",x"D6",x"03",x"B7",x"C9",x"D7", -- 0x55A0
		x"11",x"89",x"FD",x"06",x"0F",x"7E",x"A7",x"28", -- 0x55A8
		x"0D",x"FE",x"3A",x"28",x"09",x"FE",x"28",x"28", -- 0x55B0
		x"05",x"12",x"13",x"23",x"10",x"EF",x"78",x"FE", -- 0x55B8
		x"0F",x"28",x"15",x"AF",x"12",x"1B",x"1A",x"FE", -- 0x55C0
		x"20",x"28",x"F8",x"06",x"40",x"11",x"C9",x"FC", -- 0x55C8
		x"1A",x"E6",x"20",x"20",x"06",x"13",x"10",x"F8", -- 0x55D0
		x"C3",x"55",x"40",x"C5",x"D5",x"E5",x"CD",x"2A", -- 0x55D8
		x"7E",x"F5",x"4F",x"2E",x"04",x"CD",x"1A",x"7E", -- 0x55E0
		x"D5",x"DD",x"E1",x"FD",x"E1",x"E1",x"2B",x"D7", -- 0x55E8
		x"CD",x"1C",x"00",x"D1",x"C1",x"38",x"DE",x"C9", -- 0x55F0
		x"E1",x"78",x"FE",x"10",x"38",x"02",x"06",x"0F", -- 0x55F8
		x"CD",x"B7",x"7F",x"CD",x"A9",x"4E",x"12",x"23", -- 0x5600
		x"13",x"10",x"F8",x"AF",x"12",x"06",x"40",x"11", -- 0x5608
		x"C9",x"FC",x"1A",x"E6",x"40",x"20",x"06",x"13", -- 0x5610
		x"10",x"F8",x"C3",x"6B",x"6E",x"C5",x"D5",x"CD", -- 0x5618
		x"2A",x"7E",x"F5",x"4F",x"2E",x"06",x"CD",x"1A", -- 0x5620
		x"7E",x"D5",x"DD",x"E1",x"FD",x"E1",x"3E",x"FF", -- 0x5628
		x"CD",x"1C",x"00",x"D1",x"C1",x"38",x"E0",x"4F", -- 0x5630
		x"3E",x"40",x"90",x"87",x"87",x"B1",x"FE",x"09", -- 0x5638
		x"38",x"D8",x"FE",x"FC",x"30",x"D4",x"E1",x"D1", -- 0x5640
		x"A7",x"C9",x"C5",x"F5",x"1F",x"1F",x"E6",x"3F", -- 0x5648
		x"CD",x"2D",x"7E",x"F5",x"4F",x"2E",x"06",x"CD", -- 0x5650
		x"1A",x"7E",x"D5",x"DD",x"E1",x"FD",x"E1",x"F1", -- 0x5658
		x"E6",x"03",x"32",x"99",x"FD",x"C1",x"F1",x"D1", -- 0x5660
		x"E1",x"C3",x"1C",x"00",x"ED",x"53",x"56",x"F9", -- 0x5668
		x"CD",x"64",x"4C",x"E5",x"11",x"00",x"00",x"D5", -- 0x5670
		x"F5",x"CD",x"D0",x"67",x"CD",x"DF",x"2E",x"41", -- 0x5678
		x"4A",x"53",x"78",x"B1",x"28",x"06",x"7A",x"B7", -- 0x5680
		x"28",x"02",x"C5",x"D5",x"F1",x"32",x"3B",x"FB", -- 0x5688
		x"E1",x"7C",x"B5",x"20",x"0A",x"3A",x"58",x"F9", -- 0x5690
		x"B7",x"CA",x"09",x"57",x"C3",x"94",x"74",x"22", -- 0x5698
		x"3C",x"FB",x"CD",x"EE",x"56",x"28",x"E5",x"87", -- 0x56A0
		x"4F",x"2A",x"56",x"F9",x"7E",x"87",x"CC",x"5A", -- 0x56A8
		x"47",x"B9",x"28",x"05",x"23",x"23",x"23",x"18", -- 0x56B0
		x"F3",x"01",x"A2",x"56",x"C5",x"7E",x"4F",x"87", -- 0x56B8
		x"30",x"20",x"B7",x"1F",x"4F",x"C5",x"E5",x"CD", -- 0x56C0
		x"EE",x"56",x"11",x"01",x"00",x"CA",x"DF",x"56", -- 0x56C8
		x"CD",x"A8",x"64",x"D2",x"DC",x"56",x"CD",x"1C", -- 0x56D0
		x"57",x"37",x"18",x"04",x"CD",x"0B",x"57",x"B7", -- 0x56D8
		x"E1",x"C1",x"23",x"7E",x"23",x"66",x"6F",x"E9", -- 0x56E0
		x"CD",x"EE",x"56",x"28",x"C1",x"C9",x"E5",x"21", -- 0x56E8
		x"3B",x"FB",x"7E",x"B7",x"28",x"13",x"35",x"2A", -- 0x56F0
		x"3C",x"FB",x"7E",x"23",x"22",x"3C",x"FB",x"FE", -- 0x56F8
		x"20",x"28",x"EC",x"FE",x"60",x"38",x"02",x"D6", -- 0x5700
		x"20",x"E1",x"C9",x"E5",x"21",x"3B",x"FB",x"34", -- 0x5708
		x"2A",x"3C",x"FB",x"2B",x"22",x"3C",x"FB",x"E1", -- 0x5710
		x"C9",x"CD",x"E8",x"56",x"FE",x"3D",x"CA",x"7A", -- 0x5718
		x"57",x"FE",x"2B",x"28",x"F4",x"FE",x"2D",x"20", -- 0x5720
		x"06",x"11",x"95",x"57",x"D5",x"18",x"EA",x"11", -- 0x5728
		x"00",x"00",x"FE",x"2C",x"28",x"D5",x"FE",x"3B", -- 0x5730
		x"C8",x"FE",x"3A",x"30",x"CE",x"FE",x"30",x"38", -- 0x5738
		x"CA",x"21",x"00",x"00",x"06",x"0A",x"19",x"38", -- 0x5740
		x"2A",x"10",x"FB",x"D6",x"30",x"5F",x"16",x"00", -- 0x5748
		x"19",x"38",x"20",x"EB",x"CD",x"EE",x"56",x"20", -- 0x5750
		x"D9",x"C9",x"CD",x"E8",x"56",x"11",x"5E",x"F5", -- 0x5758
		x"D5",x"06",x"28",x"CD",x"A8",x"64",x"38",x"0B", -- 0x5760
		x"12",x"13",x"FE",x"3B",x"28",x"08",x"CD",x"E8", -- 0x5768
		x"56",x"10",x"F5",x"CD",x"5A",x"47",x"E1",x"C3", -- 0x5770
		x"9B",x"4E",x"CD",x"5A",x"57",x"CD",x"8A",x"2F", -- 0x5778
		x"EB",x"C9",x"CD",x"5A",x"57",x"3A",x"3B",x"FB", -- 0x5780
		x"2A",x"3C",x"FB",x"E3",x"F5",x"0E",x"02",x"CD", -- 0x5788
		x"5E",x"62",x"C3",x"79",x"56",x"AF",x"93",x"5F", -- 0x5790
		x"9A",x"93",x"57",x"C9",x"7E",x"FE",x"40",x"CC", -- 0x5798
		x"66",x"46",x"01",x"00",x"00",x"50",x"59",x"FE", -- 0x57A0
		x"F2",x"28",x"16",x"7E",x"FE",x"DC",x"F5",x"CC", -- 0x57A8
		x"66",x"46",x"CF",x"28",x"CD",x"0F",x"52",x"D5", -- 0x57B0
		x"CF",x"2C",x"CD",x"0F",x"52",x"CF",x"29",x"C1", -- 0x57B8
		x"F1",x"E5",x"2A",x"B7",x"FC",x"28",x"03",x"21", -- 0x57C0
		x"00",x"00",x"09",x"22",x"B7",x"FC",x"22",x"B3", -- 0x57C8
		x"FC",x"44",x"4D",x"2A",x"B9",x"FC",x"28",x"03", -- 0x57D0
		x"21",x"00",x"00",x"19",x"22",x"B9",x"FC",x"22", -- 0x57D8
		x"B5",x"FC",x"EB",x"E1",x"C9",x"3A",x"EA",x"F3", -- 0x57E0
		x"18",x"03",x"3A",x"E9",x"F3",x"F5",x"CD",x"AB", -- 0x57E8
		x"57",x"F1",x"CD",x"50",x"58",x"E5",x"CD",x"0E", -- 0x57F0
		x"01",x"30",x"06",x"CD",x"11",x"01",x"CD",x"20", -- 0x57F8
		x"01",x"E1",x"C9",x"D7",x"E5",x"CD",x"14",x"01", -- 0x5800
		x"D1",x"E5",x"F5",x"2A",x"B5",x"FC",x"E5",x"2A", -- 0x5808
		x"B3",x"FC",x"E5",x"2A",x"B9",x"FC",x"E5",x"2A", -- 0x5810
		x"B7",x"FC",x"E5",x"EB",x"CD",x"AB",x"57",x"E5", -- 0x5818
		x"CD",x"0E",x"01",x"21",x"FF",x"FF",x"30",x"09", -- 0x5820
		x"CD",x"11",x"01",x"CD",x"1D",x"01",x"6F",x"26", -- 0x5828
		x"00",x"CD",x"99",x"2F",x"D1",x"E1",x"22",x"B7", -- 0x5830
		x"FC",x"E1",x"22",x"B9",x"FC",x"E1",x"22",x"B3", -- 0x5838
		x"FC",x"E1",x"22",x"B5",x"FC",x"F1",x"E1",x"D5", -- 0x5840
		x"CD",x"17",x"01",x"E1",x"C9",x"3A",x"E9",x"F3", -- 0x5848
		x"C5",x"D5",x"5F",x"CD",x"BC",x"59",x"2B",x"D7", -- 0x5850
		x"28",x"09",x"CF",x"2C",x"FE",x"2C",x"28",x"03", -- 0x5858
		x"CD",x"1C",x"52",x"7B",x"E5",x"CD",x"1A",x"01", -- 0x5860
		x"DA",x"5A",x"47",x"E1",x"D1",x"C1",x"C3",x"6A", -- 0x5868
		x"46",x"2A",x"B3",x"FC",x"7D",x"91",x"6F",x"7C", -- 0x5870
		x"98",x"67",x"D0",x"AF",x"95",x"6F",x"9C",x"95", -- 0x5878
		x"67",x"37",x"C9",x"2A",x"B5",x"FC",x"7D",x"93", -- 0x5880
		x"6F",x"7C",x"9A",x"67",x"18",x"EC",x"E5",x"2A", -- 0x5888
		x"B5",x"FC",x"EB",x"22",x"B5",x"FC",x"E1",x"C9", -- 0x5890
		x"CD",x"8E",x"58",x"E5",x"C5",x"2A",x"B3",x"FC", -- 0x5898
		x"E3",x"22",x"B3",x"FC",x"C1",x"E1",x"C9",x"CD", -- 0x58A0
		x"9C",x"57",x"C5",x"D5",x"CF",x"F2",x"CD",x"AB", -- 0x58A8
		x"57",x"CD",x"4D",x"58",x"D1",x"C1",x"28",x"44", -- 0x58B0
		x"CF",x"2C",x"CF",x"42",x"CA",x"12",x"59",x"CF", -- 0x58B8
		x"46",x"E5",x"CD",x"0E",x"01",x"CD",x"98",x"58", -- 0x58C0
		x"CD",x"0E",x"01",x"CD",x"83",x"58",x"DC",x"8E", -- 0x58C8
		x"58",x"23",x"E5",x"CD",x"71",x"58",x"DC",x"9B", -- 0x58D0
		x"58",x"23",x"E5",x"CD",x"11",x"01",x"D1",x"C1", -- 0x58D8
		x"D5",x"C5",x"CD",x"14",x"01",x"F5",x"E5",x"EB", -- 0x58E0
		x"CD",x"23",x"01",x"E1",x"F1",x"CD",x"17",x"01", -- 0x58E8
		x"CD",x"08",x"01",x"C1",x"D1",x"0B",x"78",x"B1", -- 0x58F0
		x"20",x"E6",x"E1",x"C9",x"C5",x"D5",x"E5",x"CD", -- 0x58F8
		x"3C",x"59",x"2A",x"B7",x"FC",x"22",x"B3",x"FC", -- 0x5900
		x"2A",x"B9",x"FC",x"22",x"B5",x"FC",x"E1",x"D1", -- 0x5908
		x"C1",x"C9",x"E5",x"2A",x"B5",x"FC",x"E5",x"D5", -- 0x5910
		x"EB",x"CD",x"FC",x"58",x"E1",x"22",x"B5",x"FC", -- 0x5918
		x"EB",x"CD",x"FC",x"58",x"E1",x"22",x"B5",x"FC", -- 0x5920
		x"2A",x"B3",x"FC",x"C5",x"44",x"4D",x"CD",x"FC", -- 0x5928
		x"58",x"E1",x"22",x"B3",x"FC",x"44",x"4D",x"CD", -- 0x5930
		x"FC",x"58",x"E1",x"C9",x"CD",x"F3",x"FE",x"CD", -- 0x5938
		x"0E",x"01",x"CD",x"98",x"58",x"CD",x"0E",x"01", -- 0x5940
		x"CD",x"83",x"58",x"DC",x"98",x"58",x"D5",x"E5", -- 0x5948
		x"CD",x"71",x"58",x"EB",x"21",x"FC",x"00",x"30", -- 0x5950
		x"03",x"21",x"FF",x"00",x"E3",x"E7",x"30",x"10", -- 0x5958
		x"22",x"2D",x"F9",x"E1",x"22",x"ED",x"F3",x"21", -- 0x5960
		x"08",x"01",x"22",x"F0",x"F3",x"EB",x"18",x"0F", -- 0x5968
		x"E3",x"22",x"F0",x"F3",x"21",x"08",x"01",x"22", -- 0x5970
		x"ED",x"F3",x"EB",x"22",x"2D",x"F9",x"E1",x"D1", -- 0x5978
		x"E5",x"CD",x"7B",x"58",x"22",x"2F",x"F9",x"CD", -- 0x5980
		x"11",x"01",x"D1",x"D5",x"CD",x"B4",x"59",x"C1", -- 0x5988
		x"03",x"18",x"07",x"E1",x"78",x"B1",x"C8",x"CD", -- 0x5990
		x"EC",x"F3",x"CD",x"20",x"01",x"0B",x"E5",x"2A", -- 0x5998
		x"2D",x"F9",x"19",x"EB",x"2A",x"2F",x"F9",x"19", -- 0x59A0
		x"30",x"E9",x"EB",x"E1",x"78",x"B1",x"C8",x"CD", -- 0x59A8
		x"EF",x"F3",x"18",x"E3",x"7A",x"B7",x"1F",x"57", -- 0x59B0
		x"7B",x"1F",x"5F",x"C9",x"3A",x"AF",x"FC",x"FE", -- 0x59B8
		x"02",x"F0",x"C3",x"5A",x"47",x"CD",x"9C",x"57", -- 0x59C0
		x"C5",x"D5",x"CD",x"4D",x"58",x"3A",x"F2",x"F3", -- 0x59C8
		x"5F",x"2B",x"D7",x"28",x"05",x"CF",x"2C",x"CD", -- 0x59D0
		x"1C",x"52",x"7B",x"CD",x"29",x"01",x"DA",x"5A", -- 0x59D8
		x"47",x"D1",x"C1",x"E5",x"CD",x"91",x"5E",x"CD", -- 0x59E0
		x"11",x"01",x"11",x"01",x"00",x"06",x"00",x"CD", -- 0x59E8
		x"DC",x"5A",x"28",x"14",x"E5",x"CD",x"ED",x"5A", -- 0x59F0
		x"D1",x"19",x"EB",x"AF",x"CD",x"CE",x"5A",x"3E", -- 0x59F8
		x"40",x"CD",x"CE",x"5A",x"06",x"C0",x"18",x"1E", -- 0x5A00
		x"E1",x"C9",x"CD",x"BD",x"00",x"3A",x"4A",x"F9", -- 0x5A08
		x"B7",x"28",x"0C",x"2A",x"4B",x"F9",x"E5",x"2A", -- 0x5A10
		x"49",x"F9",x"E5",x"2A",x"4D",x"F9",x"E5",x"D1", -- 0x5A18
		x"C1",x"E1",x"79",x"CD",x"17",x"01",x"78",x"32", -- 0x5A20
		x"53",x"F9",x"87",x"28",x"DB",x"D5",x"30",x"05", -- 0x5A28
		x"CD",x"05",x"01",x"18",x"03",x"CD",x"0B",x"01", -- 0x5A30
		x"D1",x"38",x"E4",x"06",x"00",x"CD",x"DC",x"5A", -- 0x5A38
		x"CA",x"1F",x"5A",x"AF",x"32",x"4A",x"F9",x"CD", -- 0x5A40
		x"ED",x"5A",x"5D",x"54",x"B7",x"28",x"1A",x"2B", -- 0x5A48
		x"2B",x"7C",x"87",x"38",x"14",x"ED",x"53",x"4D", -- 0x5A50
		x"F9",x"CD",x"14",x"01",x"22",x"4B",x"F9",x"32", -- 0x5A58
		x"49",x"F9",x"3A",x"53",x"F9",x"2F",x"32",x"4A", -- 0x5A60
		x"F9",x"2A",x"51",x"F9",x"19",x"EB",x"CD",x"C2", -- 0x5A68
		x"5A",x"2A",x"42",x"F9",x"3A",x"44",x"F9",x"CD", -- 0x5A70
		x"17",x"01",x"2A",x"4F",x"F9",x"ED",x"5B",x"51", -- 0x5A78
		x"F9",x"B7",x"ED",x"52",x"28",x"39",x"38",x"1C", -- 0x5A80
		x"EB",x"06",x"01",x"CD",x"DC",x"5A",x"28",x"2F", -- 0x5A88
		x"B7",x"28",x"E7",x"EB",x"2A",x"42",x"F9",x"3A", -- 0x5A90
		x"44",x"F9",x"4F",x"3A",x"53",x"F9",x"47",x"CD", -- 0x5A98
		x"D3",x"5A",x"18",x"D6",x"CD",x"7B",x"58",x"2B", -- 0x5AA0
		x"2B",x"7C",x"87",x"38",x"12",x"23",x"E5",x"CD", -- 0x5AA8
		x"FF",x"00",x"2B",x"7C",x"B5",x"20",x"F8",x"D1", -- 0x5AB0
		x"3A",x"53",x"F9",x"2F",x"CD",x"CE",x"5A",x"C3", -- 0x5AB8
		x"0A",x"5A",x"3A",x"54",x"F9",x"4F",x"3A",x"55", -- 0x5AC0
		x"F9",x"B1",x"C8",x"3A",x"53",x"F9",x"47",x"CD", -- 0x5AC8
		x"14",x"01",x"4F",x"E3",x"C5",x"D5",x"E5",x"0E", -- 0x5AD0
		x"02",x"C3",x"5E",x"62",x"CD",x"2C",x"01",x"ED", -- 0x5AD8
		x"53",x"4F",x"F9",x"22",x"51",x"F9",x"7C",x"B5", -- 0x5AE0
		x"79",x"32",x"55",x"F9",x"C9",x"CD",x"14",x"01", -- 0x5AE8
		x"E5",x"F5",x"2A",x"42",x"F9",x"3A",x"44",x"F9", -- 0x5AF0
		x"CD",x"17",x"01",x"F1",x"E1",x"22",x"42",x"F9", -- 0x5AF8
		x"32",x"44",x"F9",x"CD",x"2F",x"01",x"79",x"32", -- 0x5B00
		x"54",x"F9",x"C9",x"EB",x"CD",x"7B",x"58",x"EB", -- 0x5B08
		x"C9",x"CD",x"9C",x"57",x"CF",x"2C",x"CD",x"0F", -- 0x5B10
		x"52",x"E5",x"EB",x"22",x"B3",x"FC",x"CD",x"99", -- 0x5B18
		x"2F",x"CD",x"B2",x"2F",x"01",x"40",x"70",x"11", -- 0x5B20
		x"71",x"07",x"CD",x"5C",x"32",x"CD",x"8A",x"2F", -- 0x5B28
		x"22",x"36",x"F9",x"AF",x"32",x"35",x"F9",x"32", -- 0x5B30
		x"41",x"F9",x"E1",x"CD",x"4D",x"58",x"0E",x"01", -- 0x5B38
		x"11",x"00",x"00",x"CD",x"17",x"5D",x"D5",x"0E", -- 0x5B40
		x"80",x"11",x"FF",x"FF",x"CD",x"17",x"5D",x"E3", -- 0x5B48
		x"AF",x"EB",x"E7",x"3E",x"00",x"30",x"0F",x"3D", -- 0x5B50
		x"EB",x"F5",x"3A",x"35",x"F9",x"4F",x"07",x"07", -- 0x5B58
		x"B1",x"0F",x"32",x"35",x"F9",x"F1",x"32",x"38", -- 0x5B60
		x"F9",x"ED",x"53",x"3F",x"F9",x"22",x"33",x"F9", -- 0x5B68
		x"E1",x"2B",x"D7",x"20",x"10",x"E5",x"CD",x"26", -- 0x5B70
		x"01",x"7C",x"B7",x"28",x"32",x"3E",x"01",x"32", -- 0x5B78
		x"41",x"F9",x"EB",x"18",x"2A",x"CF",x"2C",x"CD", -- 0x5B80
		x"64",x"4C",x"E5",x"CD",x"B2",x"2F",x"CD",x"71", -- 0x5B88
		x"2E",x"CA",x"5A",x"47",x"FA",x"5A",x"47",x"CD", -- 0x5B90
		x"63",x"5D",x"20",x"07",x"3C",x"32",x"41",x"F9", -- 0x5B98
		x"CD",x"67",x"32",x"01",x"43",x"25",x"11",x"60", -- 0x5BA0
		x"00",x"CD",x"5C",x"32",x"CD",x"8A",x"2F",x"22", -- 0x5BA8
		x"31",x"F9",x"11",x"00",x"00",x"ED",x"53",x"3D", -- 0x5BB0
		x"F9",x"2A",x"B3",x"FC",x"29",x"CD",x"BD",x"00", -- 0x5BB8
		x"7B",x"1F",x"38",x"16",x"D5",x"E5",x"23",x"EB", -- 0x5BC0
		x"CD",x"B4",x"59",x"EB",x"13",x"CD",x"B4",x"59", -- 0x5BC8
		x"CD",x"06",x"5C",x"D1",x"E1",x"E7",x"D2",x"08", -- 0x5BD0
		x"5A",x"EB",x"44",x"4D",x"2A",x"3D",x"F9",x"23", -- 0x5BD8
		x"19",x"19",x"7C",x"87",x"38",x"0C",x"D5",x"EB", -- 0x5BE0
		x"60",x"69",x"29",x"2B",x"EB",x"B7",x"ED",x"52", -- 0x5BE8
		x"0B",x"D1",x"22",x"3D",x"F9",x"60",x"69",x"13", -- 0x5BF0
		x"18",x"C3",x"D5",x"CD",x"EB",x"5C",x"E1",x"3A", -- 0x5BF8
		x"41",x"F9",x"B7",x"C8",x"EB",x"C9",x"ED",x"53", -- 0x5C00
		x"39",x"F9",x"E5",x"21",x"00",x"00",x"22",x"3B", -- 0x5C08
		x"F9",x"CD",x"FA",x"5B",x"22",x"45",x"F9",x"E1", -- 0x5C10
		x"EB",x"E5",x"CD",x"FA",x"5B",x"ED",x"53",x"47", -- 0x5C18
		x"F9",x"D1",x"CD",x"0B",x"5B",x"CD",x"48",x"5C", -- 0x5C20
		x"E5",x"D5",x"2A",x"36",x"F9",x"22",x"3B",x"F9", -- 0x5C28
		x"ED",x"5B",x"39",x"F9",x"B7",x"ED",x"52",x"22", -- 0x5C30
		x"39",x"F9",x"2A",x"45",x"F9",x"CD",x"7B",x"58", -- 0x5C38
		x"22",x"45",x"F9",x"D1",x"E1",x"CD",x"0B",x"5B", -- 0x5C40
		x"3E",x"04",x"F5",x"E5",x"D5",x"E5",x"D5",x"ED", -- 0x5C48
		x"5B",x"3B",x"F9",x"2A",x"36",x"F9",x"29",x"19", -- 0x5C50
		x"22",x"3B",x"F9",x"2A",x"39",x"F9",x"19",x"EB", -- 0x5C58
		x"2A",x"3F",x"F9",x"E7",x"28",x"1A",x"30",x"08", -- 0x5C60
		x"2A",x"33",x"F9",x"E7",x"28",x"0A",x"30",x"20", -- 0x5C68
		x"3A",x"38",x"F9",x"B7",x"20",x"24",x"18",x"1E", -- 0x5C70
		x"3A",x"35",x"F9",x"87",x"30",x"1C",x"18",x"06", -- 0x5C78
		x"3A",x"35",x"F9",x"1F",x"30",x"14",x"D1",x"E1", -- 0x5C80
		x"CD",x"DC",x"5C",x"CD",x"CD",x"5C",x"18",x"1A", -- 0x5C88
		x"3A",x"38",x"F9",x"B7",x"28",x"04",x"D1",x"E1", -- 0x5C90
		x"18",x"10",x"D1",x"E1",x"CD",x"DC",x"5C",x"CD", -- 0x5C98
		x"0E",x"01",x"30",x"06",x"CD",x"11",x"01",x"CD", -- 0x5CA0
		x"20",x"01",x"D1",x"E1",x"F1",x"3D",x"C8",x"F5", -- 0x5CA8
		x"D5",x"ED",x"5B",x"45",x"F9",x"CD",x"0B",x"5B", -- 0x5CB0
		x"22",x"45",x"F9",x"EB",x"D1",x"E5",x"2A",x"47", -- 0x5CB8
		x"F9",x"EB",x"22",x"47",x"F9",x"CD",x"0B",x"5B", -- 0x5CC0
		x"E1",x"F1",x"C3",x"4A",x"5C",x"2A",x"B7",x"FC", -- 0x5CC8
		x"22",x"B3",x"FC",x"2A",x"B9",x"FC",x"22",x"B5", -- 0x5CD0
		x"FC",x"C3",x"3C",x"59",x"D5",x"ED",x"5B",x"B7", -- 0x5CD8
		x"FC",x"19",x"44",x"4D",x"D1",x"2A",x"B9",x"FC", -- 0x5CE0
		x"19",x"EB",x"C9",x"2A",x"31",x"F9",x"7D",x"B7", -- 0x5CE8
		x"20",x"04",x"B4",x"C0",x"EB",x"C9",x"4A",x"16", -- 0x5CF0
		x"00",x"F5",x"CD",x"0A",x"5D",x"1E",x"80",x"19", -- 0x5CF8
		x"59",x"4C",x"F1",x"CD",x"0A",x"5D",x"59",x"19", -- 0x5D00
		x"EB",x"C9",x"06",x"08",x"21",x"00",x"00",x"29", -- 0x5D08
		x"87",x"30",x"01",x"19",x"10",x"F9",x"C9",x"2B", -- 0x5D10
		x"D7",x"C8",x"CF",x"2C",x"FE",x"2C",x"C8",x"C5", -- 0x5D18
		x"CD",x"64",x"4C",x"E3",x"E5",x"CD",x"B2",x"2F", -- 0x5D20
		x"C1",x"21",x"F6",x"F7",x"7E",x"B7",x"F2",x"3A", -- 0x5D28
		x"5D",x"E6",x"7F",x"77",x"21",x"35",x"F9",x"7E", -- 0x5D30
		x"B1",x"77",x"01",x"40",x"15",x"11",x"91",x"55", -- 0x5D38
		x"CD",x"5C",x"32",x"CD",x"63",x"5D",x"CA",x"5A", -- 0x5D40
		x"47",x"CD",x"B1",x"2E",x"2A",x"36",x"F9",x"29", -- 0x5D48
		x"29",x"29",x"CD",x"99",x"2F",x"CD",x"B2",x"2F", -- 0x5D50
		x"C1",x"D1",x"CD",x"5C",x"32",x"CD",x"8A",x"2F", -- 0x5D58
		x"D1",x"EB",x"C9",x"01",x"41",x"10",x"11",x"00", -- 0x5D60
		x"00",x"CD",x"21",x"2F",x"3D",x"C9",x"3A",x"AF", -- 0x5D68
		x"FC",x"FE",x"02",x"DA",x"5A",x"47",x"11",x"83", -- 0x5D70
		x"5D",x"AF",x"32",x"BB",x"FC",x"32",x"58",x"F9", -- 0x5D78
		x"C3",x"6C",x"56",x"D5",x"B1",x"5D",x"C4",x"B4", -- 0x5D80
		x"5D",x"CC",x"B9",x"5D",x"D2",x"BC",x"5D",x"4D", -- 0x5D88
		x"D8",x"5D",x"C5",x"CA",x"5D",x"C6",x"C6",x"5D", -- 0x5D90
		x"C7",x"D1",x"5D",x"C8",x"C3",x"5D",x"C1",x"4E", -- 0x5D98
		x"5E",x"42",x"46",x"5E",x"4E",x"42",x"5E",x"58", -- 0x5DA0
		x"82",x"57",x"C3",x"87",x"5E",x"D3",x"59",x"5E", -- 0x5DA8
		x"00",x"CD",x"0B",x"5B",x"01",x"00",x"00",x"18", -- 0x5DB0
		x"46",x"CD",x"0B",x"5B",x"42",x"4B",x"11",x"00", -- 0x5DB8
		x"00",x"18",x"3C",x"CD",x"0B",x"5B",x"42",x"4B", -- 0x5DC0
		x"18",x"35",x"42",x"4B",x"CD",x"0B",x"5B",x"18", -- 0x5DC8
		x"2E",x"CD",x"0B",x"5B",x"42",x"4B",x"18",x"F4", -- 0x5DD0
		x"CD",x"E8",x"56",x"06",x"00",x"FE",x"2B",x"28", -- 0x5DD8
		x"05",x"FE",x"2D",x"28",x"01",x"04",x"78",x"F5", -- 0x5DE0
		x"CD",x"0B",x"57",x"CD",x"19",x"57",x"D5",x"CD", -- 0x5DE8
		x"E8",x"56",x"FE",x"2C",x"C2",x"5A",x"47",x"CD", -- 0x5DF0
		x"19",x"57",x"C1",x"F1",x"B7",x"20",x"23",x"CD", -- 0x5DF8
		x"66",x"5E",x"D5",x"50",x"59",x"CD",x"66",x"5E", -- 0x5E00
		x"EB",x"D1",x"3A",x"BD",x"FC",x"1F",x"30",x"06", -- 0x5E08
		x"F5",x"CD",x"7B",x"58",x"EB",x"F1",x"1F",x"30", -- 0x5E10
		x"06",x"CD",x"7B",x"58",x"CD",x"0B",x"5B",x"CD", -- 0x5E18
		x"DC",x"5C",x"3A",x"BB",x"FC",x"87",x"38",x"09", -- 0x5E20
		x"F5",x"C5",x"D5",x"CD",x"CD",x"5C",x"D1",x"C1", -- 0x5E28
		x"F1",x"87",x"38",x"09",x"ED",x"53",x"B9",x"FC", -- 0x5E30
		x"60",x"69",x"22",x"B7",x"FC",x"AF",x"32",x"BB", -- 0x5E38
		x"FC",x"C9",x"3E",x"40",x"18",x"02",x"3E",x"80", -- 0x5E40
		x"21",x"BB",x"FC",x"B6",x"77",x"C9",x"30",x"09", -- 0x5E48
		x"7B",x"FE",x"04",x"30",x"04",x"32",x"BD",x"FC", -- 0x5E50
		x"C9",x"D2",x"5A",x"47",x"7A",x"B7",x"C2",x"5A", -- 0x5E58
		x"47",x"7B",x"32",x"BC",x"FC",x"C9",x"3A",x"BC", -- 0x5E60
		x"FC",x"B7",x"C8",x"21",x"00",x"00",x"19",x"3D", -- 0x5E68
		x"20",x"FC",x"EB",x"7A",x"87",x"F5",x"30",x"01", -- 0x5E70
		x"1B",x"CD",x"B4",x"59",x"CD",x"B4",x"59",x"F1", -- 0x5E78
		x"D0",x"7A",x"F6",x"C0",x"57",x"13",x"C9",x"30", -- 0x5E80
		x"D0",x"7B",x"CD",x"1A",x"01",x"DA",x"5A",x"47", -- 0x5E88
		x"C9",x"E5",x"CD",x"0E",x"01",x"D2",x"5A",x"47", -- 0x5E90
		x"E1",x"C9",x"2B",x"D7",x"C8",x"CF",x"2C",x"01", -- 0x5E98
		x"9A",x"5E",x"C5",x"F6",x"AF",x"32",x"62",x"F6", -- 0x5EA0
		x"4E",x"CD",x"A2",x"FF",x"CD",x"A7",x"64",x"DA", -- 0x5EA8
		x"55",x"40",x"AF",x"47",x"D7",x"38",x"05",x"CD", -- 0x5EB0
		x"A8",x"64",x"38",x"09",x"47",x"D7",x"38",x"FD", -- 0x5EB8
		x"CD",x"A8",x"64",x"30",x"F8",x"FE",x"26",x"30", -- 0x5EC0
		x"17",x"11",x"EE",x"5E",x"D5",x"16",x"02",x"FE", -- 0x5EC8
		x"25",x"C8",x"14",x"FE",x"24",x"C8",x"14",x"FE", -- 0x5ED0
		x"21",x"C8",x"16",x"08",x"FE",x"23",x"C8",x"F1", -- 0x5ED8
		x"79",x"E6",x"7F",x"5F",x"16",x"00",x"E5",x"21", -- 0x5EE0
		x"89",x"F6",x"19",x"56",x"E1",x"2B",x"7A",x"32", -- 0x5EE8
		x"63",x"F6",x"D7",x"3A",x"A5",x"F6",x"3D",x"CA", -- 0x5EF0
		x"E8",x"5F",x"F2",x"08",x"5F",x"7E",x"D6",x"28", -- 0x5EF8
		x"CA",x"BA",x"5F",x"D6",x"33",x"CA",x"BA",x"5F", -- 0x5F00
		x"AF",x"32",x"A5",x"F6",x"E5",x"3A",x"B7",x"F7", -- 0x5F08
		x"B7",x"32",x"B4",x"F7",x"28",x"3C",x"2A",x"E6", -- 0x5F10
		x"F6",x"11",x"E8",x"F6",x"19",x"22",x"B5",x"F7", -- 0x5F18
		x"EB",x"18",x"17",x"1A",x"6F",x"13",x"1A",x"13", -- 0x5F20
		x"B9",x"20",x"0B",x"3A",x"63",x"F6",x"BD",x"20", -- 0x5F28
		x"05",x"1A",x"B8",x"CA",x"A4",x"5F",x"13",x"26", -- 0x5F30
		x"00",x"19",x"EB",x"3A",x"B5",x"F7",x"BB",x"C2", -- 0x5F38
		x"23",x"5F",x"3A",x"B6",x"F7",x"BA",x"20",x"DB", -- 0x5F40
		x"3A",x"B4",x"F7",x"B7",x"28",x"18",x"AF",x"32", -- 0x5F48
		x"B4",x"F7",x"2A",x"C4",x"F6",x"22",x"B5",x"F7", -- 0x5F50
		x"2A",x"C2",x"F6",x"18",x"DD",x"CD",x"A4",x"5E", -- 0x5F58
		x"C9",x"57",x"5F",x"C1",x"E3",x"C9",x"E1",x"E3", -- 0x5F60
		x"D5",x"11",x"60",x"5F",x"E7",x"28",x"F2",x"11", -- 0x5F68
		x"9E",x"4E",x"E7",x"D1",x"28",x"31",x"E3",x"E5", -- 0x5F70
		x"C5",x"3A",x"63",x"F6",x"4F",x"C5",x"06",x"00", -- 0x5F78
		x"03",x"03",x"03",x"2A",x"C6",x"F6",x"E5",x"09", -- 0x5F80
		x"C1",x"E5",x"CD",x"50",x"62",x"E1",x"22",x"C6", -- 0x5F88
		x"F6",x"60",x"69",x"22",x"C4",x"F6",x"2B",x"36", -- 0x5F90
		x"00",x"E7",x"20",x"FA",x"D1",x"73",x"23",x"D1", -- 0x5F98
		x"73",x"23",x"72",x"EB",x"13",x"E1",x"C9",x"32", -- 0x5FA0
		x"F6",x"F7",x"67",x"6F",x"22",x"F8",x"F7",x"EF", -- 0x5FA8
		x"20",x"06",x"21",x"D6",x"3F",x"22",x"F8",x"F7", -- 0x5FB0
		x"E1",x"C9",x"E5",x"2A",x"62",x"F6",x"E3",x"57", -- 0x5FB8
		x"D5",x"C5",x"CD",x"55",x"47",x"C1",x"F1",x"EB", -- 0x5FC0
		x"E3",x"E5",x"EB",x"3C",x"57",x"7E",x"FE",x"2C", -- 0x5FC8
		x"CA",x"C0",x"5F",x"FE",x"29",x"28",x"05",x"FE", -- 0x5FD0
		x"5D",x"C2",x"55",x"40",x"D7",x"22",x"BC",x"F6", -- 0x5FD8
		x"E1",x"22",x"62",x"F6",x"1E",x"00",x"D5",x"11", -- 0x5FE0
		x"E5",x"F5",x"2A",x"C4",x"F6",x"3E",x"19",x"ED", -- 0x5FE8
		x"5B",x"C6",x"F6",x"E7",x"28",x"2D",x"5E",x"23", -- 0x5FF0
		x"7E",x"23",x"B9",x"20",x"08",x"3A",x"63",x"F6", -- 0x5FF8
		x"BB",x"20",x"02",x"7E",x"B8",x"23",x"5E",x"23", -- 0x6000
		x"56",x"23",x"20",x"E2",x"3A",x"62",x"F6",x"B7", -- 0x6008
		x"C2",x"5E",x"40",x"F1",x"44",x"4D",x"CA",x"97", -- 0x6010
		x"32",x"96",x"CA",x"7D",x"60",x"11",x"09",x"00", -- 0x6018
		x"C3",x"6F",x"40",x"3A",x"63",x"F6",x"77",x"23", -- 0x6020
		x"5F",x"16",x"00",x"F1",x"CA",x"5A",x"47",x"71", -- 0x6028
		x"23",x"70",x"23",x"4F",x"CD",x"5E",x"62",x"23", -- 0x6030
		x"23",x"22",x"9D",x"F6",x"71",x"23",x"3A",x"62", -- 0x6038
		x"F6",x"17",x"79",x"01",x"0B",x"00",x"30",x"02", -- 0x6040
		x"C1",x"03",x"71",x"F5",x"23",x"70",x"23",x"CD", -- 0x6048
		x"4A",x"31",x"F1",x"3D",x"20",x"ED",x"F5",x"42", -- 0x6050
		x"4B",x"EB",x"19",x"DA",x"75",x"62",x"CD",x"67", -- 0x6058
		x"62",x"22",x"C6",x"F6",x"2B",x"36",x"00",x"E7", -- 0x6060
		x"20",x"FA",x"03",x"57",x"2A",x"9D",x"F6",x"5E", -- 0x6068
		x"EB",x"29",x"09",x"EB",x"2B",x"2B",x"73",x"23", -- 0x6070
		x"72",x"23",x"F1",x"38",x"30",x"47",x"4F",x"7E", -- 0x6078
		x"23",x"16",x"E1",x"5E",x"23",x"56",x"23",x"E3", -- 0x6080
		x"F5",x"E7",x"D2",x"1D",x"60",x"CD",x"4A",x"31", -- 0x6088
		x"19",x"F1",x"3D",x"44",x"4D",x"20",x"EB",x"3A", -- 0x6090
		x"63",x"F6",x"44",x"4D",x"29",x"D6",x"04",x"38", -- 0x6098
		x"04",x"29",x"28",x"06",x"29",x"B7",x"E2",x"AA", -- 0x60A0
		x"60",x"09",x"C1",x"09",x"EB",x"2A",x"BC",x"F6", -- 0x60A8
		x"C9",x"CD",x"65",x"4C",x"CD",x"58",x"30",x"CF", -- 0x60B0
		x"3B",x"EB",x"2A",x"F8",x"F7",x"18",x"08",x"3A", -- 0x60B8
		x"A6",x"F6",x"B7",x"28",x"0D",x"D1",x"EB",x"E5", -- 0x60C0
		x"AF",x"32",x"A6",x"F6",x"3C",x"F5",x"D5",x"46", -- 0x60C8
		x"04",x"05",x"CA",x"5A",x"47",x"23",x"7E",x"23", -- 0x60D0
		x"66",x"6F",x"18",x"1A",x"58",x"E5",x"0E",x"02", -- 0x60D8
		x"7E",x"23",x"FE",x"5C",x"CA",x"10",x"62",x"FE", -- 0x60E0
		x"20",x"20",x"03",x"0C",x"10",x"F2",x"E1",x"43", -- 0x60E8
		x"3E",x"5C",x"CD",x"46",x"62",x"DF",x"AF",x"5F", -- 0x60F0
		x"57",x"CD",x"46",x"62",x"57",x"7E",x"23",x"FE", -- 0x60F8
		x"21",x"CA",x"0D",x"62",x"FE",x"23",x"28",x"3C", -- 0x6100
		x"FE",x"26",x"CA",x"09",x"62",x"05",x"CA",x"F5", -- 0x6108
		x"61",x"FE",x"2B",x"3E",x"08",x"28",x"E2",x"2B", -- 0x6110
		x"7E",x"23",x"FE",x"2E",x"28",x"40",x"FE",x"5C", -- 0x6118
		x"28",x"BA",x"BE",x"20",x"CD",x"FE",x"24",x"28", -- 0x6120
		x"14",x"FE",x"2A",x"20",x"C5",x"23",x"78",x"FE", -- 0x6128
		x"02",x"38",x"03",x"7E",x"FE",x"24",x"3E",x"20", -- 0x6130
		x"20",x"07",x"05",x"1C",x"FE",x"AF",x"C6",x"10", -- 0x6138
		x"23",x"1C",x"82",x"57",x"1C",x"0E",x"00",x"05", -- 0x6140
		x"28",x"48",x"7E",x"23",x"FE",x"2E",x"28",x"19", -- 0x6148
		x"FE",x"23",x"28",x"F0",x"FE",x"2C",x"20",x"1B", -- 0x6150
		x"7A",x"F6",x"40",x"57",x"18",x"E6",x"7E",x"FE", -- 0x6158
		x"23",x"3E",x"2E",x"C2",x"F2",x"60",x"0E",x"01", -- 0x6160
		x"23",x"0C",x"05",x"28",x"25",x"7E",x"23",x"FE", -- 0x6168
		x"23",x"28",x"F6",x"D5",x"11",x"90",x"61",x"D5", -- 0x6170
		x"54",x"5D",x"FE",x"5E",x"C0",x"BE",x"C0",x"23", -- 0x6178
		x"BE",x"C0",x"23",x"BE",x"C0",x"23",x"78",x"D6", -- 0x6180
		x"04",x"D8",x"D1",x"D1",x"47",x"14",x"23",x"CA", -- 0x6188
		x"EB",x"D1",x"7A",x"2B",x"1C",x"E6",x"08",x"20", -- 0x6190
		x"15",x"1D",x"78",x"B7",x"28",x"10",x"7E",x"D6", -- 0x6198
		x"2D",x"28",x"06",x"FE",x"FE",x"20",x"07",x"3E", -- 0x61A0
		x"08",x"C6",x"04",x"82",x"57",x"05",x"E1",x"F1", -- 0x61A8
		x"28",x"4C",x"C5",x"D5",x"CD",x"64",x"4C",x"D1", -- 0x61B0
		x"C1",x"C5",x"E5",x"43",x"78",x"81",x"FE",x"19", -- 0x61B8
		x"D2",x"5A",x"47",x"7A",x"F6",x"80",x"CD",x"26", -- 0x61C0
		x"34",x"CD",x"78",x"66",x"E1",x"2B",x"D7",x"37", -- 0x61C8
		x"28",x"0B",x"32",x"A6",x"F6",x"FE",x"3B",x"28", -- 0x61D0
		x"03",x"CF",x"2C",x"06",x"D7",x"C1",x"EB",x"E1", -- 0x61D8
		x"E5",x"F5",x"D5",x"7E",x"90",x"23",x"16",x"00", -- 0x61E0
		x"5F",x"7E",x"23",x"66",x"6F",x"19",x"78",x"B7", -- 0x61E8
		x"C2",x"F6",x"60",x"18",x"04",x"CD",x"46",x"62", -- 0x61F0
		x"DF",x"E1",x"F1",x"C2",x"BF",x"60",x"DC",x"28", -- 0x61F8
		x"73",x"E3",x"CD",x"D6",x"67",x"E1",x"C3",x"FF", -- 0x6200
		x"4A",x"0E",x"00",x"18",x"04",x"0E",x"01",x"3E", -- 0x6208
		x"F1",x"05",x"CD",x"46",x"62",x"E1",x"F1",x"28", -- 0x6210
		x"E5",x"C5",x"CD",x"64",x"4C",x"CD",x"58",x"30", -- 0x6218
		x"C1",x"C5",x"E5",x"2A",x"F8",x"F7",x"41",x"0E", -- 0x6220
		x"00",x"78",x"F5",x"B7",x"C4",x"68",x"68",x"CD", -- 0x6228
		x"7B",x"66",x"2A",x"F8",x"F7",x"F1",x"B7",x"CA", -- 0x6230
		x"CC",x"61",x"96",x"47",x"3E",x"20",x"04",x"05", -- 0x6238
		x"CA",x"CC",x"61",x"DF",x"18",x"F9",x"F5",x"7A", -- 0x6240
		x"B7",x"3E",x"2B",x"C4",x"18",x"00",x"F1",x"C9", -- 0x6248
		x"CD",x"67",x"62",x"C5",x"E3",x"C1",x"E7",x"7E", -- 0x6250
		x"02",x"C8",x"0B",x"2B",x"18",x"F8",x"E5",x"2A", -- 0x6258
		x"C6",x"F6",x"06",x"00",x"09",x"09",x"3E",x"E5", -- 0x6260
		x"3E",x"88",x"95",x"6F",x"3E",x"FF",x"9C",x"67", -- 0x6268
		x"38",x"03",x"39",x"E1",x"D8",x"CD",x"53",x"42", -- 0x6270
		x"2A",x"74",x"F6",x"2B",x"2B",x"22",x"B1",x"F6", -- 0x6278
		x"11",x"07",x"00",x"C3",x"6F",x"40",x"C0",x"2A", -- 0x6280
		x"76",x"F6",x"CD",x"39",x"64",x"32",x"AA",x"F6", -- 0x6288
		x"32",x"A9",x"F6",x"77",x"23",x"77",x"23",x"22", -- 0x6290
		x"C2",x"F6",x"CD",x"CB",x"FE",x"2A",x"76",x"F6", -- 0x6298
		x"2B",x"CD",x"D0",x"FE",x"22",x"A7",x"F6",x"CD", -- 0x62A0
		x"6E",x"63",x"06",x"1A",x"21",x"CA",x"F6",x"CD", -- 0x62A8
		x"D5",x"FE",x"36",x"08",x"23",x"10",x"FB",x"CD", -- 0x62B0
		x"24",x"2C",x"AF",x"32",x"BB",x"F6",x"6F",x"67", -- 0x62B8
		x"22",x"B9",x"F6",x"22",x"C0",x"F6",x"2A",x"72", -- 0x62C0
		x"F6",x"22",x"9B",x"F6",x"CD",x"C9",x"63",x"2A", -- 0x62C8
		x"C2",x"F6",x"22",x"C4",x"F6",x"22",x"C6",x"F6", -- 0x62D0
		x"CD",x"1C",x"6C",x"3A",x"7C",x"F8",x"E6",x"01", -- 0x62D8
		x"20",x"03",x"32",x"7C",x"F8",x"C1",x"2A",x"74", -- 0x62E0
		x"F6",x"2B",x"2B",x"22",x"B1",x"F6",x"23",x"23", -- 0x62E8
		x"CD",x"DA",x"FE",x"F9",x"21",x"7A",x"F6",x"22", -- 0x62F0
		x"78",x"F6",x"CD",x"04",x"73",x"CD",x"FF",x"4A", -- 0x62F8
		x"AF",x"67",x"6F",x"22",x"E6",x"F6",x"32",x"B7", -- 0x6300
		x"F7",x"22",x"4E",x"F7",x"22",x"BA",x"F7",x"22", -- 0x6308
		x"E4",x"F6",x"32",x"A5",x"F6",x"E5",x"C5",x"2A", -- 0x6310
		x"A7",x"F6",x"C9",x"F3",x"7E",x"E6",x"04",x"F6", -- 0x6318
		x"01",x"BE",x"77",x"28",x"04",x"E6",x"04",x"20", -- 0x6320
		x"26",x"FB",x"C9",x"F3",x"7E",x"36",x"00",x"18", -- 0x6328
		x"07",x"F3",x"7E",x"F5",x"F6",x"02",x"77",x"F1", -- 0x6330
		x"EE",x"05",x"28",x"26",x"FB",x"C9",x"F3",x"7E", -- 0x6338
		x"E6",x"05",x"BE",x"77",x"20",x"02",x"FB",x"C9", -- 0x6340
		x"EE",x"05",x"28",x"03",x"FB",x"C9",x"F3",x"3A", -- 0x6348
		x"D8",x"FB",x"3C",x"32",x"D8",x"FB",x"FB",x"C9", -- 0x6350
		x"F3",x"7E",x"E6",x"03",x"BE",x"77",x"20",x"02", -- 0x6358
		x"FB",x"C9",x"3A",x"D8",x"FB",x"D6",x"01",x"38", -- 0x6360
		x"F7",x"32",x"D8",x"FB",x"FB",x"C9",x"21",x"4C", -- 0x6368
		x"FC",x"06",x"1A",x"AF",x"77",x"23",x"77",x"23", -- 0x6370
		x"77",x"23",x"10",x"F8",x"21",x"CE",x"FB",x"06", -- 0x6378
		x"0A",x"77",x"23",x"10",x"FC",x"32",x"D8",x"FB", -- 0x6380
		x"C9",x"3A",x"BB",x"F6",x"B7",x"C0",x"E5",x"2A", -- 0x6388
		x"1C",x"F4",x"7C",x"A5",x"3C",x"28",x"0F",x"21", -- 0x6390
		x"4C",x"FC",x"06",x"1A",x"7E",x"FE",x"05",x"28", -- 0x6398
		x"07",x"23",x"23",x"23",x"10",x"F6",x"E1",x"C9", -- 0x63A0
		x"C5",x"23",x"5E",x"23",x"56",x"2B",x"2B",x"7A", -- 0x63A8
		x"B3",x"C1",x"28",x"ED",x"D5",x"E5",x"CD",x"58", -- 0x63B0
		x"63",x"CD",x"31",x"63",x"0E",x"03",x"CD",x"5E", -- 0x63B8
		x"62",x"C1",x"D1",x"E1",x"E3",x"E1",x"C3",x"CF", -- 0x63C0
		x"47",x"EB",x"2A",x"76",x"F6",x"28",x"0E",x"EB", -- 0x63C8
		x"CD",x"69",x"47",x"E5",x"CD",x"95",x"42",x"60", -- 0x63D0
		x"69",x"D1",x"D2",x"1C",x"48",x"2B",x"22",x"C8", -- 0x63D8
		x"F6",x"EB",x"C9",x"C2",x"A5",x"77",x"C0",x"3C", -- 0x63E0
		x"18",x"0A",x"C0",x"AF",x"32",x"BB",x"F6",x"F5", -- 0x63E8
		x"CC",x"1C",x"6C",x"F1",x"22",x"AF",x"F6",x"21", -- 0x63F0
		x"7A",x"F6",x"22",x"78",x"F6",x"21",x"F6",x"FF", -- 0x63F8
		x"C1",x"2A",x"1C",x"F4",x"E5",x"F5",x"7D",x"A4", -- 0x6400
		x"3C",x"28",x"09",x"22",x"BE",x"F6",x"2A",x"AF", -- 0x6408
		x"F6",x"22",x"C0",x"F6",x"CD",x"04",x"73",x"CD", -- 0x6410
		x"23",x"73",x"F1",x"21",x"DC",x"3F",x"C2",x"FD", -- 0x6418
		x"40",x"C3",x"1E",x"41",x"2A",x"C0",x"F6",x"7C", -- 0x6420
		x"B5",x"11",x"11",x"00",x"CA",x"6F",x"40",x"ED", -- 0x6428
		x"5B",x"BE",x"F6",x"ED",x"53",x"1C",x"F4",x"C9", -- 0x6430
		x"3E",x"AF",x"32",x"C4",x"F7",x"C9",x"CD",x"A4", -- 0x6438
		x"5E",x"D5",x"E5",x"21",x"BC",x"F7",x"CD",x"F3", -- 0x6440
		x"2E",x"2A",x"C4",x"F6",x"E3",x"EF",x"F5",x"CF", -- 0x6448
		x"2C",x"CD",x"A4",x"5E",x"F1",x"47",x"EF",x"B8", -- 0x6450
		x"C2",x"6D",x"40",x"E3",x"EB",x"E5",x"2A",x"C4", -- 0x6458
		x"F6",x"E7",x"20",x"10",x"D1",x"E1",x"E3",x"D5", -- 0x6460
		x"CD",x"F3",x"2E",x"E1",x"11",x"BC",x"F7",x"CD", -- 0x6468
		x"F3",x"2E",x"E1",x"C9",x"C3",x"5A",x"47",x"3E", -- 0x6470
		x"01",x"32",x"A5",x"F6",x"CD",x"A4",x"5E",x"E5", -- 0x6478
		x"32",x"A5",x"F6",x"60",x"69",x"0B",x"0B",x"0B", -- 0x6480
		x"0B",x"0B",x"19",x"EB",x"2A",x"C6",x"F6",x"E7", -- 0x6488
		x"1A",x"02",x"13",x"03",x"20",x"F9",x"0B",x"60", -- 0x6490
		x"69",x"22",x"C6",x"F6",x"E1",x"7E",x"FE",x"2C", -- 0x6498
		x"C0",x"D7",x"18",x"D3",x"F1",x"E1",x"C9",x"7E", -- 0x64A0
		x"FE",x"41",x"D8",x"FE",x"5B",x"3F",x"C9",x"CA", -- 0x64A8
		x"A1",x"62",x"CD",x"56",x"47",x"2B",x"D7",x"E5", -- 0x64B0
		x"2A",x"4A",x"FC",x"44",x"4D",x"2A",x"72",x"F6", -- 0x64B8
		x"28",x"2A",x"E1",x"CF",x"2C",x"D5",x"CD",x"2F", -- 0x64C0
		x"54",x"2B",x"D7",x"C2",x"55",x"40",x"E3",x"EB", -- 0x64C8
		x"7C",x"A7",x"F2",x"5A",x"47",x"D5",x"11",x"81", -- 0x64D0
		x"F3",x"E7",x"D2",x"5A",x"47",x"D1",x"E5",x"01", -- 0x64D8
		x"F5",x"FE",x"3A",x"5F",x"F8",x"09",x"3D",x"F2", -- 0x64E0
		x"E5",x"64",x"C1",x"2B",x"7D",x"93",x"5F",x"7C", -- 0x64E8
		x"9A",x"57",x"DA",x"75",x"62",x"E5",x"2A",x"C2", -- 0x64F0
		x"F6",x"C5",x"01",x"A0",x"00",x"09",x"C1",x"E7", -- 0x64F8
		x"D2",x"75",x"62",x"EB",x"22",x"74",x"F6",x"60", -- 0x6500
		x"69",x"22",x"4A",x"FC",x"E1",x"22",x"72",x"F6", -- 0x6508
		x"E1",x"CD",x"A1",x"62",x"3A",x"5F",x"F8",x"CD", -- 0x6510
		x"6B",x"7E",x"2A",x"A7",x"F6",x"C3",x"01",x"46", -- 0x6518
		x"7D",x"93",x"5F",x"7C",x"9A",x"57",x"C9",x"11", -- 0x6520
		x"00",x"00",x"C4",x"A4",x"5E",x"22",x"A7",x"F6", -- 0x6528
		x"CD",x"E2",x"3F",x"C2",x"5B",x"40",x"F9",x"D5", -- 0x6530
		x"7E",x"F5",x"23",x"D5",x"7E",x"23",x"B7",x"FA", -- 0x6538
		x"6B",x"65",x"3D",x"20",x"04",x"01",x"08",x"00", -- 0x6540
		x"09",x"C6",x"04",x"32",x"63",x"F6",x"CD",x"08", -- 0x6548
		x"2F",x"EB",x"E3",x"E5",x"EF",x"30",x"4E",x"CD", -- 0x6550
		x"D6",x"2E",x"CD",x"4E",x"32",x"E1",x"CD",x"E8", -- 0x6558
		x"2E",x"E1",x"CD",x"DF",x"2E",x"E5",x"CD",x"21", -- 0x6560
		x"2F",x"18",x"29",x"01",x"0C",x"00",x"09",x"4E", -- 0x6568
		x"23",x"46",x"23",x"E3",x"5E",x"23",x"56",x"E5", -- 0x6570
		x"69",x"60",x"CD",x"72",x"31",x"3A",x"63",x"F6", -- 0x6578
		x"FE",x"02",x"C2",x"67",x"40",x"EB",x"E1",x"72", -- 0x6580
		x"2B",x"73",x"E1",x"D5",x"5E",x"23",x"56",x"23", -- 0x6588
		x"E3",x"CD",x"4D",x"2F",x"E1",x"C1",x"90",x"CD", -- 0x6590
		x"DF",x"2E",x"28",x"1A",x"EB",x"22",x"1C",x"F4", -- 0x6598
		x"69",x"60",x"C3",x"FD",x"45",x"CD",x"97",x"26", -- 0x65A0
		x"E1",x"CD",x"10",x"2F",x"E1",x"CD",x"EF",x"2E", -- 0x65A8
		x"D5",x"CD",x"5C",x"2F",x"18",x"DE",x"F9",x"22", -- 0x65B0
		x"B1",x"F6",x"EB",x"2A",x"A7",x"F6",x"7E",x"FE", -- 0x65B8
		x"2C",x"C2",x"01",x"46",x"D7",x"CD",x"2A",x"65", -- 0x65C0
		x"CD",x"D0",x"67",x"7E",x"23",x"4E",x"23",x"46", -- 0x65C8
		x"D1",x"C5",x"F5",x"CD",x"D7",x"67",x"F1",x"57", -- 0x65D0
		x"5E",x"23",x"4E",x"23",x"46",x"E1",x"7B",x"B2", -- 0x65D8
		x"C8",x"7A",x"D6",x"01",x"D8",x"AF",x"BB",x"3C", -- 0x65E0
		x"D0",x"15",x"1D",x"0A",x"03",x"BE",x"23",x"28", -- 0x65E8
		x"ED",x"3F",x"C3",x"79",x"2E",x"CD",x"1E",x"37", -- 0x65F0
		x"18",x"0D",x"CD",x"22",x"37",x"18",x"08",x"CD", -- 0x65F8
		x"1A",x"37",x"18",x"03",x"CD",x"25",x"34",x"CD", -- 0x6600
		x"35",x"66",x"CD",x"D3",x"67",x"01",x"25",x"68", -- 0x6608
		x"C5",x"7E",x"23",x"E5",x"CD",x"8E",x"66",x"E1", -- 0x6610
		x"4E",x"23",x"46",x"CD",x"2A",x"66",x"E5",x"6F", -- 0x6618
		x"CD",x"C7",x"67",x"D1",x"C9",x"3E",x"01",x"CD", -- 0x6620
		x"8E",x"66",x"21",x"98",x"F6",x"E5",x"77",x"23", -- 0x6628
		x"73",x"23",x"72",x"E1",x"C9",x"2B",x"06",x"22", -- 0x6630
		x"50",x"E5",x"0E",x"FF",x"23",x"7E",x"0C",x"B7", -- 0x6638
		x"28",x"06",x"BA",x"28",x"03",x"B8",x"20",x"F4", -- 0x6640
		x"FE",x"22",x"CC",x"66",x"46",x"E3",x"23",x"EB", -- 0x6648
		x"79",x"CD",x"2A",x"66",x"11",x"98",x"F6",x"3E", -- 0x6650
		x"D5",x"2A",x"78",x"F6",x"22",x"F8",x"F7",x"3E", -- 0x6658
		x"03",x"32",x"63",x"F6",x"CD",x"F3",x"2E",x"11", -- 0x6660
		x"9B",x"F6",x"E7",x"22",x"78",x"F6",x"E1",x"7E", -- 0x6668
		x"C0",x"11",x"10",x"00",x"C3",x"6F",x"40",x"23", -- 0x6670
		x"CD",x"35",x"66",x"CD",x"D3",x"67",x"CD",x"E1", -- 0x6678
		x"2E",x"14",x"15",x"C8",x"0A",x"DF",x"FE",x"0D", -- 0x6680
		x"CC",x"31",x"73",x"03",x"18",x"F4",x"B7",x"0E", -- 0x6688
		x"F1",x"F5",x"2A",x"74",x"F6",x"EB",x"2A",x"9B", -- 0x6690
		x"F6",x"2F",x"4F",x"06",x"FF",x"09",x"23",x"E7", -- 0x6698
		x"38",x"07",x"22",x"9B",x"F6",x"23",x"EB",x"F1", -- 0x66A0
		x"C9",x"F1",x"11",x"0E",x"00",x"CA",x"6F",x"40", -- 0x66A8
		x"BF",x"F5",x"01",x"90",x"66",x"C5",x"2A",x"72", -- 0x66B0
		x"F6",x"22",x"9B",x"F6",x"21",x"00",x"00",x"E5", -- 0x66B8
		x"2A",x"C6",x"F6",x"E5",x"21",x"7A",x"F6",x"ED", -- 0x66C0
		x"5B",x"78",x"F6",x"E7",x"01",x"C7",x"66",x"C2", -- 0x66C8
		x"42",x"67",x"21",x"4C",x"F7",x"22",x"B8",x"F7", -- 0x66D0
		x"2A",x"C4",x"F6",x"22",x"B5",x"F7",x"2A",x"C2", -- 0x66D8
		x"F6",x"ED",x"5B",x"B5",x"F7",x"E7",x"28",x"12", -- 0x66E0
		x"7E",x"23",x"23",x"23",x"FE",x"03",x"20",x"04", -- 0x66E8
		x"CD",x"43",x"67",x"AF",x"5F",x"16",x"00",x"19", -- 0x66F0
		x"18",x"E7",x"2A",x"B8",x"F7",x"5E",x"23",x"56", -- 0x66F8
		x"7A",x"B3",x"2A",x"C4",x"F6",x"28",x"13",x"EB", -- 0x6700
		x"22",x"B8",x"F7",x"23",x"23",x"5E",x"23",x"56", -- 0x6708
		x"23",x"EB",x"19",x"22",x"B5",x"F7",x"EB",x"18", -- 0x6710
		x"C8",x"C1",x"ED",x"5B",x"C6",x"F6",x"E7",x"CA", -- 0x6718
		x"63",x"67",x"7E",x"23",x"CD",x"DF",x"2E",x"E5", -- 0x6720
		x"09",x"FE",x"03",x"20",x"EC",x"22",x"9F",x"F6", -- 0x6728
		x"E1",x"4E",x"06",x"00",x"09",x"09",x"23",x"EB", -- 0x6730
		x"2A",x"9F",x"F6",x"EB",x"E7",x"28",x"DB",x"01", -- 0x6738
		x"37",x"67",x"C5",x"AF",x"B6",x"23",x"5E",x"23", -- 0x6740
		x"56",x"23",x"C8",x"44",x"4D",x"2A",x"9B",x"F6", -- 0x6748
		x"E7",x"60",x"69",x"D8",x"E1",x"E3",x"E7",x"E3", -- 0x6750
		x"E5",x"60",x"69",x"D0",x"C1",x"F1",x"F1",x"E5", -- 0x6758
		x"D5",x"C5",x"C9",x"D1",x"E1",x"7C",x"B5",x"C8", -- 0x6760
		x"2B",x"46",x"2B",x"4E",x"E5",x"2B",x"6E",x"26", -- 0x6768
		x"00",x"09",x"50",x"59",x"2B",x"44",x"4D",x"2A", -- 0x6770
		x"9B",x"F6",x"CD",x"53",x"62",x"E1",x"71",x"23", -- 0x6778
		x"70",x"60",x"69",x"2B",x"C3",x"B9",x"66",x"C5", -- 0x6780
		x"E5",x"2A",x"F8",x"F7",x"E3",x"CD",x"C7",x"4D", -- 0x6788
		x"E3",x"CD",x"58",x"30",x"7E",x"E5",x"2A",x"F8", -- 0x6790
		x"F7",x"E5",x"86",x"11",x"0F",x"00",x"DA",x"6F", -- 0x6798
		x"40",x"CD",x"27",x"66",x"D1",x"CD",x"D7",x"67", -- 0x67A0
		x"E3",x"CD",x"D6",x"67",x"E5",x"2A",x"99",x"F6", -- 0x67A8
		x"EB",x"CD",x"BF",x"67",x"CD",x"BF",x"67",x"21", -- 0x67B0
		x"73",x"4C",x"E3",x"E5",x"C3",x"54",x"66",x"E1", -- 0x67B8
		x"E3",x"7E",x"23",x"4E",x"23",x"46",x"6F",x"2C", -- 0x67C0
		x"2D",x"C8",x"0A",x"12",x"03",x"13",x"18",x"F8", -- 0x67C8
		x"CD",x"58",x"30",x"2A",x"F8",x"F7",x"EB",x"CD", -- 0x67D0
		x"EE",x"67",x"EB",x"C0",x"D5",x"50",x"59",x"1B", -- 0x67D8
		x"4E",x"2A",x"9B",x"F6",x"E7",x"20",x"05",x"47", -- 0x67E0
		x"09",x"22",x"9B",x"F6",x"E1",x"C9",x"CD",x"9D", -- 0x67E8
		x"FF",x"2A",x"78",x"F6",x"2B",x"46",x"2B",x"4E", -- 0x67F0
		x"2B",x"E7",x"C0",x"22",x"78",x"F6",x"C9",x"01", -- 0x67F8
		x"CF",x"4F",x"C5",x"CD",x"D0",x"67",x"AF",x"57", -- 0x6800
		x"7E",x"B7",x"C9",x"01",x"CF",x"4F",x"C5",x"CD", -- 0x6808
		x"03",x"68",x"CA",x"5A",x"47",x"23",x"5E",x"23", -- 0x6810
		x"56",x"1A",x"C9",x"CD",x"25",x"66",x"CD",x"1F", -- 0x6818
		x"52",x"2A",x"99",x"F6",x"73",x"C1",x"C3",x"54", -- 0x6820
		x"66",x"D7",x"CF",x"28",x"CD",x"1C",x"52",x"D5", -- 0x6828
		x"CF",x"2C",x"CD",x"64",x"4C",x"CF",x"29",x"E3", -- 0x6830
		x"E5",x"EF",x"28",x"05",x"CD",x"1F",x"52",x"18", -- 0x6838
		x"03",x"CD",x"0F",x"68",x"D1",x"CD",x"4D",x"68", -- 0x6840
		x"CD",x"1F",x"52",x"3E",x"20",x"F5",x"7B",x"CD", -- 0x6848
		x"27",x"66",x"47",x"F1",x"04",x"05",x"28",x"CD", -- 0x6850
		x"2A",x"99",x"F6",x"77",x"23",x"10",x"FC",x"18", -- 0x6858
		x"C4",x"CD",x"E3",x"68",x"AF",x"E3",x"4F",x"3E", -- 0x6860
		x"E5",x"E5",x"7E",x"B8",x"38",x"02",x"78",x"11", -- 0x6868
		x"0E",x"00",x"C5",x"CD",x"8E",x"66",x"C1",x"E1", -- 0x6870
		x"E5",x"23",x"46",x"23",x"66",x"68",x"06",x"00", -- 0x6878
		x"09",x"44",x"4D",x"CD",x"2A",x"66",x"6F",x"CD", -- 0x6880
		x"C7",x"67",x"D1",x"CD",x"D7",x"67",x"C3",x"54", -- 0x6888
		x"66",x"CD",x"E3",x"68",x"D1",x"D5",x"1A",x"90", -- 0x6890
		x"18",x"CB",x"EB",x"7E",x"CD",x"E6",x"68",x"04", -- 0x6898
		x"05",x"CA",x"5A",x"47",x"C5",x"CD",x"E4",x"69", -- 0x68A0
		x"F1",x"E3",x"01",x"69",x"68",x"C5",x"3D",x"BE", -- 0x68A8
		x"06",x"00",x"D0",x"4F",x"7E",x"91",x"BB",x"47", -- 0x68B0
		x"D8",x"43",x"C9",x"CD",x"03",x"68",x"CA",x"CF", -- 0x68B8
		x"4F",x"5F",x"23",x"7E",x"23",x"66",x"6F",x"E5", -- 0x68C0
		x"19",x"46",x"22",x"19",x"F4",x"78",x"32",x"1B", -- 0x68C8
		x"F4",x"72",x"E3",x"C5",x"2B",x"D7",x"CD",x"99", -- 0x68D0
		x"32",x"21",x"00",x"00",x"22",x"19",x"F4",x"C1", -- 0x68D8
		x"E1",x"70",x"C9",x"EB",x"CF",x"29",x"C1",x"D1", -- 0x68E0
		x"C5",x"43",x"C9",x"D7",x"CD",x"62",x"4C",x"EF", -- 0x68E8
		x"3E",x"01",x"F5",x"28",x"11",x"F1",x"CD",x"1F", -- 0x68F0
		x"52",x"B7",x"CA",x"5A",x"47",x"F5",x"CF",x"2C", -- 0x68F8
		x"CD",x"64",x"4C",x"CD",x"58",x"30",x"CF",x"2C", -- 0x6900
		x"E5",x"2A",x"F8",x"F7",x"E3",x"CD",x"64",x"4C", -- 0x6908
		x"CF",x"29",x"E5",x"CD",x"D0",x"67",x"EB",x"C1", -- 0x6910
		x"E1",x"F1",x"C5",x"01",x"97",x"32",x"C5",x"01", -- 0x6918
		x"CF",x"4F",x"C5",x"F5",x"D5",x"CD",x"D6",x"67", -- 0x6920
		x"D1",x"F1",x"47",x"3D",x"4F",x"BE",x"3E",x"00", -- 0x6928
		x"D0",x"1A",x"B7",x"78",x"C8",x"7E",x"23",x"46", -- 0x6930
		x"23",x"66",x"68",x"06",x"00",x"09",x"91",x"47", -- 0x6938
		x"C5",x"D5",x"E3",x"4E",x"23",x"5E",x"23",x"56", -- 0x6940
		x"E1",x"E5",x"D5",x"C5",x"1A",x"BE",x"20",x"16", -- 0x6948
		x"13",x"0D",x"28",x"09",x"23",x"10",x"F5",x"D1", -- 0x6950
		x"D1",x"C1",x"D1",x"AF",x"C9",x"E1",x"D1",x"D1", -- 0x6958
		x"C1",x"78",x"94",x"81",x"3C",x"C9",x"C1",x"D1", -- 0x6960
		x"E1",x"23",x"10",x"DD",x"18",x"EC",x"CF",x"28", -- 0x6968
		x"CD",x"A4",x"5E",x"CD",x"58",x"30",x"E5",x"D5", -- 0x6970
		x"EB",x"23",x"5E",x"23",x"56",x"2A",x"C6",x"F6", -- 0x6978
		x"E7",x"38",x"10",x"2A",x"76",x"F6",x"E7",x"30", -- 0x6980
		x"0A",x"E1",x"E5",x"CD",x"11",x"66",x"E1",x"E5", -- 0x6988
		x"CD",x"F3",x"2E",x"E1",x"E3",x"CF",x"2C",x"CD", -- 0x6990
		x"1C",x"52",x"B7",x"CA",x"5A",x"47",x"F5",x"7E", -- 0x6998
		x"CD",x"E4",x"69",x"D5",x"CD",x"5F",x"4C",x"E5", -- 0x69A0
		x"CD",x"D0",x"67",x"EB",x"E1",x"C1",x"F1",x"47", -- 0x69A8
		x"E3",x"E5",x"21",x"97",x"32",x"E3",x"79",x"B7", -- 0x69B0
		x"C8",x"7E",x"90",x"DA",x"5A",x"47",x"3C",x"B9", -- 0x69B8
		x"38",x"01",x"79",x"48",x"0D",x"06",x"00",x"D5", -- 0x69C0
		x"23",x"5E",x"23",x"66",x"6B",x"09",x"47",x"D1", -- 0x69C8
		x"EB",x"4E",x"23",x"7E",x"23",x"66",x"6F",x"EB", -- 0x69D0
		x"79",x"B7",x"C8",x"1A",x"77",x"13",x"23",x"0D", -- 0x69D8
		x"C8",x"10",x"F8",x"C9",x"1E",x"FF",x"FE",x"29", -- 0x69E0
		x"28",x"05",x"CF",x"2C",x"CD",x"1C",x"52",x"CF", -- 0x69E8
		x"29",x"C9",x"2A",x"C6",x"F6",x"EB",x"21",x"00", -- 0x69F0
		x"00",x"39",x"EF",x"C2",x"C1",x"4F",x"CD",x"D3", -- 0x69F8
		x"67",x"CD",x"B6",x"66",x"ED",x"5B",x"74",x"F6", -- 0x6A00
		x"2A",x"9B",x"F6",x"C3",x"C1",x"4F",x"CD",x"64", -- 0x6A08
		x"4C",x"E5",x"CD",x"D0",x"67",x"7E",x"B7",x"28", -- 0x6A10
		x"2E",x"23",x"5E",x"23",x"66",x"6B",x"5F",x"CD", -- 0x6A18
		x"15",x"6F",x"F5",x"01",x"66",x"F8",x"16",x"0B", -- 0x6A20
		x"1C",x"1D",x"28",x"35",x"7E",x"FE",x"20",x"38", -- 0x6A28
		x"16",x"FE",x"2E",x"28",x"18",x"02",x"03",x"23", -- 0x6A30
		x"15",x"20",x"EE",x"F1",x"F5",x"57",x"3A",x"66", -- 0x6A38
		x"F8",x"3C",x"28",x"03",x"F1",x"E1",x"C9",x"C3", -- 0x6A40
		x"6B",x"6E",x"23",x"18",x"DC",x"7A",x"FE",x"0B", -- 0x6A48
		x"CA",x"47",x"6A",x"FE",x"03",x"DA",x"47",x"6A", -- 0x6A50
		x"28",x"F0",x"3E",x"20",x"02",x"03",x"15",x"18", -- 0x6A58
		x"EC",x"3E",x"20",x"02",x"03",x"15",x"20",x"F9", -- 0x6A60
		x"18",x"D1",x"CD",x"1F",x"52",x"6F",x"3A",x"5F", -- 0x6A68
		x"F8",x"BD",x"DA",x"7D",x"6E",x"26",x"00",x"29", -- 0x6A70
		x"EB",x"2A",x"60",x"F8",x"19",x"7E",x"23",x"66", -- 0x6A78
		x"6F",x"3A",x"7C",x"F8",x"3C",x"C8",x"7E",x"B7", -- 0x6A80
		x"C8",x"E5",x"11",x"04",x"00",x"19",x"7E",x"FE", -- 0x6A88
		x"09",x"30",x"06",x"CD",x"4E",x"FE",x"C3",x"80", -- 0x6A90
		x"6E",x"E1",x"7E",x"B7",x"37",x"C9",x"2B",x"D7", -- 0x6A98
		x"FE",x"23",x"CC",x"66",x"46",x"CD",x"1C",x"52", -- 0x6AA0
		x"E3",x"E5",x"CD",x"6D",x"6A",x"CA",x"77",x"6E", -- 0x6AA8
		x"22",x"64",x"F8",x"CD",x"53",x"FE",x"C9",x"01", -- 0x6AB0
		x"FF",x"4A",x"C5",x"CD",x"0E",x"6A",x"7E",x"FE", -- 0x6AB8
		x"82",x"1E",x"04",x"20",x"1F",x"D7",x"FE",x"85", -- 0x6AC0
		x"1E",x"01",x"28",x"17",x"FE",x"9C",x"28",x"0C", -- 0x6AC8
		x"CF",x"41",x"CF",x"50",x"CF",x"50",x"CF",x"81", -- 0x6AD0
		x"1E",x"08",x"18",x"08",x"D7",x"CF",x"B3",x"1E", -- 0x6AD8
		x"02",x"18",x"01",x"D7",x"CF",x"41",x"CF",x"53", -- 0x6AE0
		x"D5",x"7E",x"FE",x"23",x"CC",x"66",x"46",x"CD", -- 0x6AE8
		x"1C",x"52",x"B7",x"CA",x"7D",x"6E",x"CD",x"58", -- 0x6AF0
		x"FE",x"1E",x"D5",x"2B",x"5F",x"D7",x"C2",x"55", -- 0x6AF8
		x"40",x"E3",x"7B",x"F5",x"E5",x"CD",x"6D",x"6A", -- 0x6B00
		x"C2",x"6E",x"6E",x"D1",x"7A",x"FE",x"09",x"CD", -- 0x6B08
		x"5D",x"FE",x"DA",x"80",x"6E",x"E5",x"01",x"04", -- 0x6B10
		x"00",x"09",x"72",x"3E",x"00",x"E1",x"CD",x"8F", -- 0x6B18
		x"6F",x"F1",x"E1",x"C9",x"E5",x"B7",x"20",x"08", -- 0x6B20
		x"3A",x"7C",x"F8",x"E6",x"01",x"C2",x"F3",x"6C", -- 0x6B28
		x"CD",x"6D",x"6A",x"28",x"15",x"22",x"64",x"F8", -- 0x6B30
		x"E5",x"38",x"06",x"CD",x"62",x"FE",x"C3",x"80", -- 0x6B38
		x"6E",x"3E",x"02",x"CD",x"8F",x"6F",x"CD",x"EA", -- 0x6B40
		x"6C",x"E1",x"E5",x"11",x"07",x"00",x"19",x"77", -- 0x6B48
		x"67",x"6F",x"22",x"64",x"F8",x"E1",x"86",x"36", -- 0x6B50
		x"00",x"E1",x"C9",x"37",x"11",x"F6",x"AF",x"F5", -- 0x6B58
		x"CD",x"0E",x"6A",x"CD",x"67",x"FE",x"F1",x"F5", -- 0x6B60
		x"28",x"0C",x"7E",x"D6",x"2C",x"B7",x"20",x"06", -- 0x6B68
		x"D7",x"CF",x"52",x"F1",x"37",x"F5",x"F5",x"AF", -- 0x6B70
		x"1E",x"01",x"CD",x"FA",x"6A",x"2A",x"64",x"F8", -- 0x6B78
		x"01",x"07",x"00",x"09",x"F1",x"9F",x"E6",x"80", -- 0x6B80
		x"F6",x"01",x"32",x"7C",x"F8",x"F1",x"F5",x"9F", -- 0x6B88
		x"32",x"66",x"F8",x"7E",x"B7",x"FA",x"D4",x"6B", -- 0x6B90
		x"F1",x"C4",x"87",x"62",x"AF",x"CD",x"AA",x"6A", -- 0x6B98
		x"C3",x"34",x"41",x"CD",x"0E",x"6A",x"CD",x"6C", -- 0x6BA0
		x"FE",x"2B",x"D7",x"1E",x"80",x"37",x"28",x"07", -- 0x6BA8
		x"CF",x"2C",x"CF",x"41",x"B7",x"1E",x"02",x"F5", -- 0x6BB0
		x"7A",x"FE",x"09",x"38",x"05",x"1E",x"02",x"F1", -- 0x6BB8
		x"AF",x"F5",x"AF",x"CD",x"FA",x"6A",x"F1",x"38", -- 0x6BC0
		x"05",x"2B",x"D7",x"C3",x"2E",x"52",x"CD",x"71", -- 0x6BC8
		x"FE",x"C3",x"6B",x"6E",x"CD",x"76",x"FE",x"C3", -- 0x6BD0
		x"6B",x"6E",x"E5",x"D5",x"2A",x"64",x"F8",x"11", -- 0x6BD8
		x"04",x"00",x"19",x"7E",x"D1",x"E1",x"C9",x"20", -- 0x6BE0
		x"19",x"E5",x"C5",x"F5",x"11",x"F3",x"6B",x"D5", -- 0x6BE8
		x"C5",x"B7",x"C9",x"F1",x"C1",x"3D",x"F2",x"EA", -- 0x6BF0
		x"6B",x"E1",x"C9",x"C1",x"E1",x"7E",x"FE",x"2C", -- 0x6BF8
		x"C0",x"D7",x"C5",x"7E",x"FE",x"23",x"CC",x"66", -- 0x6C00
		x"46",x"CD",x"1C",x"52",x"E3",x"E5",x"11",x"FB", -- 0x6C08
		x"6B",x"D5",x"37",x"E9",x"01",x"24",x"6B",x"3A", -- 0x6C10
		x"5F",x"F8",x"18",x"CB",x"3A",x"7C",x"F8",x"B7", -- 0x6C18
		x"F8",x"01",x"24",x"6B",x"AF",x"3A",x"5F",x"F8", -- 0x6C20
		x"18",x"BD",x"3E",x"01",x"32",x"16",x"F4",x"CD", -- 0x6C28
		x"7B",x"FE",x"C3",x"5A",x"47",x"F5",x"CD",x"9E", -- 0x6C30
		x"6A",x"38",x"06",x"CD",x"80",x"FE",x"C3",x"6B", -- 0x6C38
		x"6E",x"D1",x"C1",x"3E",x"04",x"C3",x"8F",x"6F", -- 0x6C40
		x"E5",x"D5",x"C5",x"F5",x"CD",x"62",x"6C",x"30", -- 0x6C48
		x"06",x"CD",x"85",x"FE",x"C3",x"6B",x"6E",x"F1", -- 0x6C50
		x"F5",x"4F",x"3E",x"06",x"CD",x"8F",x"6F",x"C3", -- 0x6C58
		x"FF",x"72",x"D5",x"2A",x"64",x"F8",x"EB",x"21", -- 0x6C60
		x"04",x"00",x"19",x"7E",x"EB",x"D1",x"FE",x"09", -- 0x6C68
		x"C9",x"E5",x"D5",x"C5",x"CD",x"62",x"6C",x"30", -- 0x6C70
		x"06",x"CD",x"8A",x"FE",x"C3",x"80",x"6E",x"3E", -- 0x6C78
		x"08",x"CD",x"8F",x"6F",x"C3",x"00",x"73",x"D7", -- 0x6C80
		x"CF",x"24",x"CF",x"28",x"E5",x"2A",x"64",x"F8", -- 0x6C88
		x"E5",x"21",x"00",x"00",x"22",x"64",x"F8",x"E1", -- 0x6C90
		x"E3",x"CD",x"1C",x"52",x"D5",x"7E",x"FE",x"2C", -- 0x6C98
		x"20",x"11",x"D7",x"CD",x"9E",x"6A",x"FE",x"01", -- 0x6CA0
		x"CA",x"B0",x"6C",x"FE",x"04",x"C2",x"83",x"6E", -- 0x6CA8
		x"E1",x"AF",x"7E",x"F5",x"CF",x"29",x"F1",x"E3", -- 0x6CB0
		x"F5",x"7D",x"B7",x"CA",x"5A",x"47",x"E5",x"CD", -- 0x6CB8
		x"27",x"66",x"EB",x"C1",x"F1",x"F5",x"28",x"1A", -- 0x6CC0
		x"CD",x"9F",x"00",x"F5",x"CD",x"BD",x"00",x"F1", -- 0x6CC8
		x"77",x"23",x"0D",x"20",x"EF",x"F1",x"C1",x"E1", -- 0x6CD0
		x"CD",x"8F",x"FE",x"22",x"64",x"F8",x"C5",x"C3", -- 0x6CD8
		x"54",x"66",x"CD",x"71",x"6C",x"DA",x"83",x"6E", -- 0x6CE0
		x"18",x"E6",x"CD",x"FB",x"6C",x"E5",x"06",x"00", -- 0x6CE8
		x"CD",x"F5",x"6C",x"E1",x"C9",x"AF",x"77",x"23", -- 0x6CF0
		x"10",x"FC",x"C9",x"2A",x"64",x"F8",x"11",x"09", -- 0x6CF8
		x"00",x"19",x"C9",x"CD",x"94",x"FE",x"CD",x"6A", -- 0x6D00
		x"6A",x"28",x"20",x"3E",x"0A",x"38",x"21",x"CD", -- 0x6D08
		x"99",x"FE",x"18",x"22",x"CD",x"94",x"FE",x"CD", -- 0x6D10
		x"6A",x"6A",x"28",x"0F",x"3E",x"0C",x"38",x"10", -- 0x6D18
		x"CD",x"9E",x"FE",x"18",x"11",x"CD",x"94",x"FE", -- 0x6D20
		x"CD",x"6A",x"6A",x"CA",x"77",x"6E",x"3E",x"0E", -- 0x6D28
		x"DA",x"8F",x"6F",x"CD",x"A3",x"FE",x"C3",x"80", -- 0x6D30
		x"6E",x"CD",x"94",x"FE",x"CD",x"6A",x"6A",x"3E", -- 0x6D38
		x"10",x"38",x"ED",x"CD",x"A8",x"FE",x"18",x"EE", -- 0x6D40
		x"CD",x"4A",x"01",x"CA",x"40",x"46",x"AF",x"CD", -- 0x6D48
		x"24",x"6B",x"C3",x"71",x"6E",x"0E",x"01",x"FE", -- 0x6D50
		x"23",x"C0",x"C5",x"CD",x"1B",x"52",x"CF",x"2C", -- 0x6D58
		x"7B",x"E5",x"CD",x"AA",x"6A",x"7E",x"E1",x"C1", -- 0x6D60
		x"B9",x"28",x"0E",x"FE",x"04",x"28",x"0A",x"FE", -- 0x6D68
		x"08",x"20",x"03",x"79",x"FE",x"02",x"C2",x"7D", -- 0x6D70
		x"6E",x"7E",x"C9",x"01",x"17",x"63",x"C5",x"AF", -- 0x6D78
		x"C3",x"24",x"6B",x"EF",x"01",x"F1",x"4B",x"11", -- 0x6D80
		x"20",x"2C",x"20",x"17",x"5A",x"18",x"14",x"01", -- 0x6D88
		x"FF",x"4A",x"C5",x"CD",x"55",x"6D",x"CD",x"A4", -- 0x6D90
		x"5E",x"CD",x"58",x"30",x"D5",x"01",x"7B",x"48", -- 0x6D98
		x"AF",x"57",x"5F",x"F5",x"C5",x"E5",x"CD",x"71", -- 0x6DA0
		x"6C",x"DA",x"83",x"6E",x"FE",x"20",x"20",x"04", -- 0x6DA8
		x"14",x"15",x"20",x"F2",x"FE",x"22",x"20",x"0E", -- 0x6DB0
		x"7B",x"FE",x"2C",x"3E",x"22",x"20",x"07",x"57", -- 0x6DB8
		x"5F",x"CD",x"71",x"6C",x"38",x"47",x"21",x"5E", -- 0x6DC0
		x"F5",x"06",x"FF",x"4F",x"7A",x"FE",x"22",x"79", -- 0x6DC8
		x"28",x"2A",x"FE",x"0D",x"E5",x"28",x"50",x"E1", -- 0x6DD0
		x"FE",x"0A",x"20",x"20",x"4F",x"7B",x"FE",x"2C", -- 0x6DD8
		x"79",x"C4",x"61",x"6E",x"CD",x"71",x"6C",x"38", -- 0x6DE0
		x"24",x"FE",x"0A",x"28",x"EF",x"FE",x"0D",x"20", -- 0x6DE8
		x"0B",x"7B",x"FE",x"20",x"28",x"12",x"FE",x"2C", -- 0x6DF0
		x"3E",x"0D",x"28",x"0C",x"B7",x"28",x"09",x"BA", -- 0x6DF8
		x"28",x"0B",x"BB",x"28",x"08",x"CD",x"61",x"6E", -- 0x6E00
		x"CD",x"71",x"6C",x"30",x"BE",x"E5",x"FE",x"22", -- 0x6E08
		x"28",x"04",x"FE",x"20",x"20",x"2B",x"CD",x"71", -- 0x6E10
		x"6C",x"38",x"26",x"FE",x"20",x"28",x"F7",x"FE", -- 0x6E18
		x"2C",x"28",x"1E",x"FE",x"0D",x"20",x"09",x"CD", -- 0x6E20
		x"71",x"6C",x"38",x"15",x"FE",x"0A",x"28",x"11", -- 0x6E28
		x"4F",x"CD",x"62",x"6C",x"30",x"06",x"CD",x"AD", -- 0x6E30
		x"FE",x"C3",x"80",x"6E",x"3E",x"12",x"CD",x"8F", -- 0x6E38
		x"6F",x"E1",x"36",x"00",x"21",x"5D",x"F5",x"7B", -- 0x6E40
		x"D6",x"20",x"28",x"07",x"06",x"00",x"CD",x"38", -- 0x6E48
		x"66",x"E1",x"C9",x"EF",x"F5",x"D7",x"F1",x"F5", -- 0x6E50
		x"DC",x"99",x"32",x"F1",x"D4",x"99",x"32",x"E1", -- 0x6E58
		x"C9",x"B7",x"C8",x"77",x"23",x"05",x"C0",x"F1", -- 0x6E60
		x"C3",x"42",x"6E",x"1E",x"38",x"01",x"1E",x"36", -- 0x6E68
		x"01",x"1E",x"39",x"01",x"1E",x"35",x"01",x"1E", -- 0x6E70
		x"3B",x"01",x"1E",x"32",x"01",x"1E",x"34",x"01", -- 0x6E78
		x"1E",x"33",x"01",x"1E",x"37",x"01",x"1E",x"3A", -- 0x6E80
		x"AF",x"32",x"7C",x"F8",x"32",x"AE",x"FC",x"C3", -- 0x6E88
		x"6F",x"40",x"CD",x"0E",x"6A",x"D5",x"CF",x"2C", -- 0x6E90
		x"CD",x"0B",x"6F",x"EB",x"22",x"BF",x"FC",x"EB", -- 0x6E98
		x"D5",x"CF",x"2C",x"CD",x"0B",x"6F",x"EB",x"22", -- 0x6EA0
		x"7D",x"F8",x"EB",x"2B",x"D7",x"28",x"0A",x"CF", -- 0x6EA8
		x"2C",x"CD",x"0B",x"6F",x"EB",x"22",x"BF",x"FC", -- 0x6EB0
		x"EB",x"C1",x"D1",x"E5",x"C5",x"7A",x"FE",x"FF", -- 0x6EB8
		x"CA",x"D7",x"6F",x"C3",x"6B",x"6E",x"CD",x"0E", -- 0x6EC0
		x"6A",x"D5",x"AF",x"32",x"BE",x"FC",x"2B",x"D7", -- 0x6EC8
		x"01",x"00",x"00",x"28",x"13",x"CF",x"2C",x"FE", -- 0x6ED0
		x"52",x"20",x"08",x"32",x"BE",x"FC",x"D7",x"28", -- 0x6ED8
		x"07",x"CF",x"2C",x"CD",x"0B",x"6F",x"42",x"4B", -- 0x6EE0
		x"D1",x"E5",x"C5",x"7A",x"FE",x"FF",x"CA",x"14", -- 0x6EE8
		x"70",x"C3",x"6B",x"6E",x"3A",x"BE",x"FC",x"B7", -- 0x6EF0
		x"28",x"0C",x"AF",x"CD",x"24",x"6B",x"21",x"F3", -- 0x6EF8
		x"6C",x"E5",x"2A",x"BF",x"FC",x"E9",x"E1",x"AF", -- 0x6F00
		x"C3",x"24",x"6B",x"CD",x"64",x"4C",x"E5",x"CD", -- 0x6F08
		x"39",x"54",x"D1",x"EB",x"C9",x"CD",x"B2",x"FE", -- 0x6F10
		x"7E",x"FE",x"3A",x"38",x"1A",x"E5",x"53",x"7E", -- 0x6F18
		x"23",x"1D",x"28",x"0A",x"FE",x"3A",x"28",x"15", -- 0x6F20
		x"7E",x"23",x"1D",x"F2",x"24",x"6F",x"5A",x"E1", -- 0x6F28
		x"AF",x"3E",x"FF",x"CD",x"B7",x"FE",x"C9",x"CD", -- 0x6F30
		x"BC",x"FE",x"C3",x"6B",x"6E",x"7A",x"93",x"3D", -- 0x6F38
		x"C1",x"D5",x"C5",x"4F",x"47",x"11",x"76",x"6F", -- 0x6F40
		x"E3",x"E5",x"CD",x"A9",x"4E",x"C5",x"47",x"1A", -- 0x6F48
		x"23",x"13",x"B8",x"C1",x"20",x"0D",x"0D",x"20", -- 0x6F50
		x"F1",x"1A",x"B7",x"F2",x"63",x"6F",x"E1",x"E1", -- 0x6F58
		x"D1",x"B7",x"C9",x"B7",x"FA",x"59",x"6F",x"1A", -- 0x6F60
		x"87",x"13",x"30",x"FB",x"48",x"E1",x"E5",x"1A", -- 0x6F68
		x"B7",x"20",x"D7",x"C3",x"F8",x"55",x"43",x"41", -- 0x6F70
		x"53",x"FF",x"4C",x"50",x"54",x"FE",x"43",x"52", -- 0x6F78
		x"54",x"FD",x"47",x"52",x"50",x"FC",x"00",x"C7", -- 0x6F80
		x"71",x"A6",x"72",x"A2",x"71",x"82",x"71",x"CD", -- 0x6F88
		x"C6",x"FE",x"E5",x"D5",x"F5",x"11",x"04",x"00", -- 0x6F90
		x"19",x"7E",x"FE",x"FC",x"DA",x"4A",x"56",x"3E", -- 0x6F98
		x"FF",x"96",x"87",x"5F",x"21",x"87",x"6F",x"19", -- 0x6FA0
		x"5E",x"23",x"56",x"F1",x"6F",x"26",x"00",x"19", -- 0x6FA8
		x"5E",x"23",x"56",x"EB",x"D1",x"E3",x"C9",x"CD", -- 0x6FB0
		x"98",x"70",x"2B",x"D7",x"28",x"05",x"CF",x"2C", -- 0x6FB8
		x"CD",x"2D",x"7A",x"E5",x"3E",x"D3",x"CD",x"25", -- 0x6FC0
		x"71",x"2A",x"C2",x"F6",x"22",x"7D",x"F8",x"2A", -- 0x6FC8
		x"76",x"F6",x"CD",x"3E",x"71",x"E1",x"C9",x"3E", -- 0x6FD0
		x"D0",x"CD",x"25",x"71",x"AF",x"CD",x"F8",x"72", -- 0x6FD8
		x"E1",x"E5",x"CD",x"03",x"70",x"2A",x"7D",x"F8", -- 0x6FE0
		x"E5",x"CD",x"03",x"70",x"2A",x"BF",x"FC",x"CD", -- 0x6FE8
		x"03",x"70",x"D1",x"E1",x"7E",x"CD",x"DE",x"72", -- 0x6FF0
		x"E7",x"30",x"03",x"23",x"18",x"F6",x"CD",x"F0", -- 0x6FF8
		x"00",x"E1",x"C9",x"7D",x"CD",x"DE",x"72",x"7C", -- 0x7000
		x"C3",x"DE",x"72",x"CD",x"D4",x"72",x"6F",x"CD", -- 0x7008
		x"D4",x"72",x"67",x"C9",x"0E",x"D0",x"CD",x"B8", -- 0x7010
		x"70",x"CD",x"E9",x"72",x"C1",x"CD",x"0B",x"70", -- 0x7018
		x"09",x"EB",x"CD",x"0B",x"70",x"09",x"E5",x"CD", -- 0x7020
		x"0B",x"70",x"22",x"BF",x"FC",x"EB",x"D1",x"CD", -- 0x7028
		x"D4",x"72",x"77",x"E7",x"28",x"03",x"23",x"18", -- 0x7030
		x"F6",x"CD",x"E7",x"00",x"C3",x"F4",x"6E",x"D6", -- 0x7038
		x"91",x"28",x"02",x"AF",x"01",x"2F",x"23",x"FE", -- 0x7040
		x"01",x"F5",x"CD",x"8C",x"70",x"0E",x"D3",x"CD", -- 0x7048
		x"B8",x"70",x"F1",x"32",x"F8",x"F7",x"DC",x"87", -- 0x7050
		x"62",x"3A",x"F8",x"F7",x"FE",x"01",x"32",x"F5", -- 0x7058
		x"F3",x"F5",x"CD",x"EA",x"54",x"F1",x"2A",x"76", -- 0x7060
		x"F6",x"CD",x"5D",x"71",x"20",x"10",x"22",x"C2", -- 0x7068
		x"F6",x"21",x"D7",x"3F",x"CD",x"78",x"66",x"2A", -- 0x7070
		x"76",x"F6",x"E5",x"C3",x"37",x"42",x"23",x"EB", -- 0x7078
		x"2A",x"C2",x"F6",x"E7",x"DA",x"71",x"70",x"1E", -- 0x7080
		x"14",x"C3",x"6F",x"40",x"2B",x"D7",x"20",x"08", -- 0x7088
		x"E5",x"21",x"66",x"F8",x"06",x"06",x"18",x"19", -- 0x7090
		x"CD",x"64",x"4C",x"E5",x"CD",x"0F",x"68",x"2B", -- 0x7098
		x"2B",x"46",x"0E",x"06",x"21",x"66",x"F8",x"1A", -- 0x70A0
		x"77",x"23",x"13",x"0D",x"28",x"08",x"10",x"F7", -- 0x70A8
		x"41",x"36",x"20",x"23",x"10",x"FB",x"E1",x"C9", -- 0x70B0
		x"CD",x"E9",x"72",x"06",x"0A",x"CD",x"D4",x"72", -- 0x70B8
		x"B9",x"20",x"F5",x"10",x"F8",x"21",x"71",x"F8", -- 0x70C0
		x"E5",x"06",x"06",x"CD",x"D4",x"72",x"77",x"23", -- 0x70C8
		x"10",x"F9",x"E1",x"11",x"66",x"F8",x"06",x"06", -- 0x70D0
		x"1A",x"13",x"FE",x"20",x"20",x"04",x"10",x"F8", -- 0x70D8
		x"18",x"0D",x"11",x"66",x"F8",x"06",x"06",x"1A", -- 0x70E0
		x"BE",x"20",x"0A",x"23",x"13",x"10",x"F8",x"21", -- 0x70E8
		x"FF",x"70",x"C3",x"0D",x"71",x"C5",x"21",x"06", -- 0x70F0
		x"71",x"CD",x"0D",x"71",x"C1",x"18",x"B9",x"46", -- 0x70F8
		x"6F",x"75",x"6E",x"64",x"3A",x"00",x"53",x"6B", -- 0x7100
		x"69",x"70",x"20",x"3A",x"00",x"ED",x"5B",x"1C", -- 0x7108
		x"F4",x"13",x"7A",x"B3",x"C0",x"CD",x"78",x"66", -- 0x7110
		x"21",x"71",x"F8",x"06",x"06",x"7E",x"23",x"DF", -- 0x7118
		x"10",x"FB",x"C3",x"28",x"73",x"CD",x"F8",x"72", -- 0x7120
		x"06",x"0A",x"CD",x"DE",x"72",x"10",x"FB",x"06", -- 0x7128
		x"06",x"21",x"66",x"F8",x"7E",x"23",x"CD",x"DE", -- 0x7130
		x"72",x"10",x"F9",x"C3",x"F0",x"00",x"E5",x"CD", -- 0x7138
		x"EA",x"54",x"AF",x"CD",x"F8",x"72",x"D1",x"2A", -- 0x7140
		x"7D",x"F8",x"1A",x"13",x"CD",x"DE",x"72",x"E7", -- 0x7148
		x"20",x"F8",x"2E",x"07",x"CD",x"DE",x"72",x"2D", -- 0x7150
		x"20",x"FA",x"C3",x"F0",x"00",x"CD",x"E9",x"72", -- 0x7158
		x"9F",x"2F",x"57",x"06",x"0A",x"CD",x"D4",x"72", -- 0x7160
		x"5F",x"CD",x"67",x"62",x"7B",x"96",x"A2",x"C2", -- 0x7168
		x"E7",x"00",x"73",x"7E",x"B7",x"23",x"20",x"EB", -- 0x7170
		x"10",x"EB",x"01",x"FA",x"FF",x"09",x"AF",x"C3", -- 0x7178
		x"E7",x"00",x"B6",x"71",x"C2",x"71",x"86",x"6E", -- 0x7180
		x"96",x"71",x"5A",x"47",x"5A",x"47",x"5A",x"47", -- 0x7188
		x"5A",x"47",x"5A",x"47",x"5A",x"47",x"3A",x"AF", -- 0x7190
		x"FC",x"FE",x"02",x"DA",x"5A",x"47",x"79",x"C3", -- 0x7198
		x"8D",x"00",x"B6",x"71",x"C2",x"71",x"86",x"6E", -- 0x71A0
		x"C3",x"71",x"5A",x"47",x"5A",x"47",x"5A",x"47", -- 0x71A8
		x"5A",x"47",x"5A",x"47",x"5A",x"47",x"CD",x"CD", -- 0x71B0
		x"72",x"FE",x"01",x"CA",x"6B",x"6E",x"22",x"64", -- 0x71B8
		x"F8",x"73",x"C9",x"79",x"C3",x"A2",x"00",x"DB", -- 0x71C0
		x"71",x"05",x"72",x"86",x"6E",x"2A",x"72",x"3F", -- 0x71C8
		x"72",x"5A",x"47",x"5A",x"47",x"6D",x"72",x"5A", -- 0x71D0
		x"47",x"7C",x"72",x"E5",x"D5",x"01",x"06",x"00", -- 0x71D8
		x"09",x"AF",x"77",x"32",x"B1",x"FC",x"CD",x"CD", -- 0x71E0
		x"72",x"FE",x"04",x"CA",x"6B",x"6E",x"FE",x"01", -- 0x71E8
		x"28",x"09",x"3E",x"EA",x"CD",x"25",x"71",x"D1", -- 0x71F0
		x"E1",x"18",x"C3",x"0E",x"EA",x"CD",x"B8",x"70", -- 0x71F8
		x"CD",x"E7",x"00",x"18",x"F2",x"7E",x"FE",x"01", -- 0x7200
		x"28",x"1B",x"3E",x"1A",x"E5",x"CD",x"8B",x"72", -- 0x7208
		x"CC",x"2F",x"72",x"E1",x"CD",x"81",x"72",x"28", -- 0x7210
		x"0C",x"E5",x"09",x"36",x"1A",x"23",x"0C",x"20", -- 0x7218
		x"FA",x"E1",x"CD",x"2F",x"72",x"AF",x"32",x"B1", -- 0x7220
		x"FC",x"C9",x"79",x"CD",x"8B",x"72",x"C0",x"AF", -- 0x7228
		x"CD",x"F8",x"72",x"06",x"00",x"7E",x"CD",x"DE", -- 0x7230
		x"72",x"23",x"10",x"F9",x"C3",x"F0",x"00",x"EB", -- 0x7238
		x"21",x"B1",x"FC",x"CD",x"BE",x"72",x"EB",x"CD", -- 0x7240
		x"9B",x"72",x"20",x"14",x"E5",x"CD",x"E9",x"72", -- 0x7248
		x"E1",x"06",x"00",x"CD",x"D4",x"72",x"77",x"23", -- 0x7250
		x"10",x"F9",x"CD",x"E7",x"00",x"25",x"AF",x"47", -- 0x7258
		x"4F",x"09",x"7E",x"FE",x"1A",x"37",x"3F",x"C0", -- 0x7260
		x"32",x"B1",x"FC",x"37",x"C9",x"CD",x"3F",x"72", -- 0x7268
		x"21",x"B1",x"FC",x"77",x"D6",x"1A",x"D6",x"01", -- 0x7270
		x"9F",x"C3",x"9A",x"2E",x"21",x"B1",x"FC",x"71", -- 0x7278
		x"C9",x"01",x"06",x"00",x"09",x"7E",x"4F",x"36", -- 0x7280
		x"00",x"18",x"16",x"5F",x"01",x"06",x"00",x"09", -- 0x7288
		x"7E",x"34",x"23",x"23",x"23",x"E5",x"4F",x"09", -- 0x7290
		x"73",x"E1",x"C9",x"01",x"06",x"00",x"09",x"7E", -- 0x7298
		x"34",x"23",x"23",x"23",x"A7",x"C9",x"B6",x"71", -- 0x72A0
		x"C2",x"71",x"86",x"6E",x"BA",x"72",x"5A",x"47", -- 0x72A8
		x"5A",x"47",x"5A",x"47",x"5A",x"47",x"5A",x"47", -- 0x72B0
		x"5A",x"47",x"79",x"C3",x"4D",x"01",x"7E",x"36", -- 0x72B8
		x"00",x"A7",x"C8",x"33",x"33",x"FE",x"1A",x"37", -- 0x72C0
		x"3F",x"C0",x"77",x"37",x"C9",x"7B",x"FE",x"08", -- 0x72C8
		x"CA",x"6B",x"6E",x"C9",x"E5",x"D5",x"C5",x"CD", -- 0x72D0
		x"E4",x"00",x"30",x"24",x"18",x"14",x"E5",x"D5", -- 0x72D8
		x"C5",x"F5",x"CD",x"ED",x"00",x"30",x"18",x"18", -- 0x72E0
		x"09",x"E5",x"D5",x"C5",x"F5",x"CD",x"E1",x"00", -- 0x72E8
		x"30",x"0D",x"CD",x"E7",x"00",x"C3",x"B2",x"73", -- 0x72F0
		x"E5",x"D5",x"C5",x"F5",x"CD",x"EA",x"00",x"F1", -- 0x72F8
		x"C1",x"D1",x"E1",x"C9",x"AF",x"32",x"16",x"F4", -- 0x7300
		x"3A",x"15",x"F4",x"B7",x"C8",x"3E",x"0D",x"CD", -- 0x7308
		x"1C",x"73",x"3E",x"0A",x"CD",x"1C",x"73",x"AF", -- 0x7310
		x"32",x"15",x"F4",x"C9",x"CD",x"A5",x"00",x"D0", -- 0x7318
		x"C3",x"B2",x"73",x"3A",x"61",x"F6",x"B7",x"C8", -- 0x7320
		x"CD",x"E9",x"FE",x"3E",x"0D",x"DF",x"3E",x"0A", -- 0x7328
		x"DF",x"CD",x"4A",x"01",x"28",x"02",x"AF",x"C9", -- 0x7330
		x"3A",x"16",x"F4",x"B7",x"28",x"05",x"AF",x"32", -- 0x7338
		x"15",x"F4",x"C9",x"32",x"61",x"F6",x"C9",x"D7", -- 0x7340
		x"E5",x"CD",x"9C",x"00",x"28",x"0C",x"CD",x"9F", -- 0x7348
		x"00",x"F5",x"CD",x"25",x"66",x"F1",x"5F",x"CD", -- 0x7350
		x"21",x"68",x"21",x"D6",x"3F",x"22",x"F8",x"F7", -- 0x7358
		x"3E",x"03",x"32",x"63",x"F6",x"E1",x"C9",x"DF", -- 0x7360
		x"FE",x"0A",x"C0",x"3E",x"0D",x"DF",x"CD",x"31", -- 0x7368
		x"73",x"3E",x"0A",x"C9",x"CD",x"EE",x"FE",x"06", -- 0x7370
		x"FF",x"21",x"5E",x"F5",x"CD",x"71",x"6C",x"38", -- 0x7378
		x"16",x"77",x"FE",x"0D",x"28",x"0B",x"FE",x"09", -- 0x7380
		x"28",x"04",x"FE",x"0A",x"28",x"EE",x"23",x"10", -- 0x7388
		x"EB",x"AF",x"77",x"21",x"5D",x"F5",x"C9",x"04", -- 0x7390
		x"20",x"F7",x"3A",x"7C",x"F8",x"E6",x"80",x"32", -- 0x7398
		x"7C",x"F8",x"CD",x"7B",x"6D",x"3A",x"66",x"F8", -- 0x73A0
		x"A7",x"CA",x"1E",x"41",x"CD",x"9A",x"62",x"C3", -- 0x73A8
		x"01",x"46",x"1E",x"13",x"C3",x"6F",x"40",x"1E", -- 0x73B0
		x"FF",x"28",x"0B",x"D6",x"EB",x"5F",x"28",x"05", -- 0x73B8
		x"CF",x"95",x"1E",x"01",x"3E",x"D7",x"7B",x"C3", -- 0x73C0
		x"F3",x"00",x"CD",x"1C",x"52",x"FE",x"0E",x"D2", -- 0x73C8
		x"5A",x"47",x"F5",x"CF",x"2C",x"CD",x"1C",x"52", -- 0x73D0
		x"F1",x"FE",x"07",x"20",x"04",x"CB",x"B3",x"CB", -- 0x73D8
		x"FB",x"C3",x"93",x"00",x"20",x"CD",x"C5",x"FF", -- 0x73E0
		x"E5",x"21",x"2E",x"75",x"22",x"56",x"F9",x"3E", -- 0x73E8
		x"00",x"32",x"35",x"FB",x"21",x"F6",x"FF",x"39", -- 0x73F0
		x"22",x"36",x"FB",x"E1",x"F5",x"CD",x"64",x"4C", -- 0x73F8
		x"E3",x"E5",x"CD",x"D0",x"67",x"CD",x"DF",x"2E", -- 0x7400
		x"7B",x"B7",x"20",x"07",x"1E",x"01",x"01",x"E4", -- 0x7408
		x"73",x"51",x"48",x"F1",x"F5",x"CD",x"50",x"01", -- 0x7410
		x"73",x"23",x"72",x"23",x"71",x"23",x"54",x"5D", -- 0x7418
		x"01",x"1C",x"00",x"09",x"EB",x"73",x"23",x"72", -- 0x7420
		x"C1",x"E1",x"04",x"78",x"FE",x"03",x"30",x"16", -- 0x7428
		x"2B",x"D7",x"28",x"05",x"C5",x"CF",x"2C",x"18", -- 0x7430
		x"C4",x"78",x"32",x"38",x"FB",x"CD",x"07",x"75", -- 0x7438
		x"04",x"78",x"FE",x"03",x"38",x"F3",x"2B",x"D7", -- 0x7440
		x"C2",x"55",x"40",x"E5",x"AF",x"F5",x"32",x"38", -- 0x7448
		x"FB",x"47",x"CD",x"21",x"75",x"DA",x"D6",x"74", -- 0x7450
		x"78",x"CD",x"50",x"01",x"7E",x"B7",x"CA",x"D6", -- 0x7458
		x"74",x"32",x"3B",x"FB",x"23",x"5E",x"23",x"56", -- 0x7460
		x"23",x"ED",x"53",x"3C",x"FB",x"5E",x"23",x"56", -- 0x7468
		x"23",x"E5",x"2E",x"24",x"CD",x"53",x"01",x"E5", -- 0x7470
		x"2A",x"36",x"FB",x"2B",x"C1",x"F3",x"CD",x"53", -- 0x7478
		x"62",x"D1",x"60",x"69",x"F9",x"FB",x"3E",x"FF", -- 0x7480
		x"32",x"58",x"F9",x"C3",x"A2",x"56",x"3A",x"3B", -- 0x7488
		x"FB",x"B7",x"20",x"03",x"CD",x"07",x"75",x"3A", -- 0x7490
		x"38",x"FB",x"CD",x"50",x"01",x"3A",x"3B",x"FB", -- 0x7498
		x"77",x"23",x"ED",x"5B",x"3C",x"FB",x"73",x"23", -- 0x74A0
		x"72",x"21",x"00",x"00",x"39",x"EB",x"2A",x"36", -- 0x74A8
		x"FB",x"F3",x"F9",x"C1",x"C1",x"C1",x"E5",x"B7", -- 0x74B0
		x"ED",x"52",x"28",x"18",x"3E",x"F0",x"A5",x"B4", -- 0x74B8
		x"C2",x"5A",x"47",x"2E",x"24",x"CD",x"53",x"01", -- 0x74C0
		x"C1",x"0B",x"CD",x"53",x"62",x"E1",x"2B",x"70", -- 0x74C8
		x"2B",x"71",x"18",x"02",x"C1",x"C1",x"FB",x"F1", -- 0x74D0
		x"3C",x"FE",x"03",x"DA",x"4D",x"74",x"F3",x"3A", -- 0x74D8
		x"9B",x"FC",x"FE",x"03",x"28",x"1C",x"3A",x"35", -- 0x74E0
		x"FB",x"07",x"38",x"07",x"21",x"40",x"FB",x"34", -- 0x74E8
		x"CD",x"99",x"00",x"FB",x"21",x"35",x"FB",x"7E", -- 0x74F0
		x"F6",x"80",x"77",x"FE",x"83",x"C2",x"4C",x"74", -- 0x74F8
		x"E1",x"C9",x"CD",x"90",x"00",x"18",x"F9",x"3A", -- 0x7500
		x"35",x"FB",x"3C",x"32",x"35",x"FB",x"1E",x"FF", -- 0x7508
		x"E5",x"C5",x"D5",x"3A",x"38",x"FB",x"F3",x"CD", -- 0x7510
		x"F9",x"00",x"FB",x"D1",x"28",x"F4",x"C1",x"E1", -- 0x7518
		x"C9",x"3A",x"38",x"FB",x"C5",x"F3",x"CD",x"F6", -- 0x7520
		x"00",x"FB",x"C1",x"FE",x"08",x"C9",x"41",x"3E", -- 0x7528
		x"76",x"42",x"3E",x"76",x"43",x"3E",x"76",x"44", -- 0x7530
		x"3E",x"76",x"45",x"3E",x"76",x"46",x"3E",x"76", -- 0x7538
		x"47",x"3E",x"76",x"CD",x"9E",x"75",x"D6",x"86", -- 0x7540
		x"75",x"D3",x"BE",x"75",x"CE",x"21",x"76",x"CF", -- 0x7548
		x"EF",x"75",x"D2",x"FC",x"75",x"D4",x"E2",x"75", -- 0x7550
		x"CC",x"C8",x"75",x"58",x"82",x"57",x"00",x"10", -- 0x7558
		x"12",x"14",x"16",x"00",x"00",x"02",x"04",x"06", -- 0x7560
		x"08",x"0A",x"0A",x"0C",x"0E",x"10",x"5D",x"0D", -- 0x7568
		x"9C",x"0C",x"E7",x"0B",x"3C",x"0B",x"9B",x"0A", -- 0x7570
		x"02",x"0A",x"73",x"09",x"EB",x"08",x"6B",x"08", -- 0x7578
		x"F2",x"07",x"80",x"07",x"14",x"07",x"38",x"02", -- 0x7580
		x"1E",x"08",x"3E",x"0F",x"BB",x"38",x"50",x"AF", -- 0x7588
		x"B2",x"20",x"4C",x"2E",x"12",x"CD",x"53",x"01", -- 0x7590
		x"3E",x"40",x"A6",x"B3",x"77",x"C9",x"7B",x"38", -- 0x7598
		x"03",x"2F",x"3C",x"5F",x"B2",x"28",x"38",x"2E", -- 0x75A0
		x"13",x"CD",x"53",x"01",x"E5",x"7E",x"23",x"66", -- 0x75A8
		x"6F",x"E7",x"E1",x"C8",x"73",x"23",x"72",x"2B", -- 0x75B0
		x"2B",x"3E",x"40",x"B6",x"77",x"C9",x"7B",x"FE", -- 0x75B8
		x"10",x"30",x"1C",x"F6",x"10",x"5F",x"18",x"C7", -- 0x75C0
		x"38",x"02",x"1E",x"04",x"7B",x"FE",x"41",x"30", -- 0x75C8
		x"0E",x"2E",x"10",x"CD",x"53",x"01",x"AF",x"B2", -- 0x75D0
		x"20",x"05",x"B3",x"28",x"02",x"77",x"C9",x"CD", -- 0x75D8
		x"5A",x"47",x"38",x"02",x"1E",x"78",x"7B",x"FE", -- 0x75E0
		x"20",x"38",x"F4",x"2E",x"11",x"18",x"E4",x"38", -- 0x75E8
		x"02",x"1E",x"04",x"7B",x"FE",x"09",x"30",x"E7", -- 0x75F0
		x"2E",x"0F",x"18",x"D7",x"38",x"02",x"1E",x"04", -- 0x75F8
		x"AF",x"B2",x"20",x"DB",x"B3",x"28",x"D8",x"FE", -- 0x7600
		x"41",x"30",x"D4",x"21",x"00",x"00",x"E5",x"2E", -- 0x7608
		x"10",x"CD",x"53",x"01",x"E5",x"23",x"23",x"7E", -- 0x7610
		x"32",x"39",x"FB",x"36",x"80",x"2B",x"2B",x"18", -- 0x7618
		x"7B",x"30",x"BC",x"AF",x"B2",x"20",x"B8",x"B3", -- 0x7620
		x"28",x"E1",x"FE",x"61",x"30",x"B1",x"7B",x"06", -- 0x7628
		x"00",x"58",x"D6",x"0C",x"1C",x"30",x"FB",x"C6", -- 0x7630
		x"0C",x"87",x"4F",x"C3",x"73",x"76",x"41",x"79", -- 0x7638
		x"D6",x"40",x"87",x"4F",x"CD",x"EE",x"56",x"28", -- 0x7640
		x"1C",x"FE",x"23",x"28",x"19",x"FE",x"2B",x"28", -- 0x7648
		x"15",x"FE",x"2D",x"28",x"05",x"CD",x"0B",x"57", -- 0x7650
		x"18",x"0B",x"0D",x"78",x"FE",x"43",x"28",x"04", -- 0x7658
		x"FE",x"46",x"20",x"01",x"0D",x"0D",x"2E",x"0F", -- 0x7660
		x"CD",x"53",x"01",x"5E",x"06",x"00",x"21",x"5F", -- 0x7668
		x"75",x"09",x"4E",x"21",x"6E",x"75",x"09",x"7B", -- 0x7670
		x"5E",x"23",x"56",x"3D",x"28",x"09",x"CB",x"3A", -- 0x7678
		x"CB",x"1B",x"18",x"F7",x"CD",x"5A",x"47",x"8B", -- 0x7680
		x"5F",x"8A",x"93",x"57",x"D5",x"2E",x"10",x"CD", -- 0x7688
		x"53",x"01",x"4E",x"E5",x"CD",x"EE",x"56",x"28", -- 0x7690
		x"10",x"CD",x"2F",x"57",x"3E",x"40",x"BB",x"38", -- 0x7698
		x"E3",x"AF",x"B2",x"20",x"DF",x"B3",x"28",x"01", -- 0x76A0
		x"4B",x"E1",x"16",x"00",x"42",x"23",x"5E",x"E5", -- 0x76A8
		x"CD",x"4A",x"31",x"EB",x"CD",x"CB",x"2F",x"CD", -- 0x76B0
		x"0D",x"2F",x"21",x"54",x"77",x"CD",x"BE",x"2E", -- 0x76B8
		x"CD",x"9F",x"28",x"CD",x"8A",x"2F",x"54",x"5D", -- 0x76C0
		x"CD",x"EE",x"56",x"28",x"16",x"FE",x"2E",x"20", -- 0x76C8
		x"0F",x"CB",x"3A",x"CB",x"1B",x"ED",x"5A",x"3E", -- 0x76D0
		x"E0",x"A4",x"28",x"EC",x"AC",x"67",x"18",x"03", -- 0x76D8
		x"CD",x"0B",x"57",x"11",x"05",x"00",x"E7",x"38", -- 0x76E0
		x"01",x"EB",x"01",x"F7",x"FF",x"E1",x"E5",x"09", -- 0x76E8
		x"72",x"23",x"73",x"23",x"0E",x"02",x"E3",x"23", -- 0x76F0
		x"5E",x"7B",x"E6",x"BF",x"77",x"E3",x"3E",x"80", -- 0x76F8
		x"B3",x"77",x"23",x"0C",x"E3",x"7B",x"E6",x"40", -- 0x7700
		x"28",x"0C",x"23",x"5E",x"23",x"56",x"E1",x"72", -- 0x7708
		x"23",x"73",x"23",x"0C",x"0C",x"FE",x"E1",x"D1", -- 0x7710
		x"7A",x"B3",x"28",x"05",x"72",x"23",x"73",x"0C", -- 0x7718
		x"0C",x"2E",x"07",x"CD",x"53",x"01",x"71",x"79", -- 0x7720
		x"D6",x"02",x"0F",x"0F",x"0F",x"23",x"B6",x"77", -- 0x7728
		x"2B",x"7A",x"B3",x"20",x"0C",x"E5",x"3A",x"39", -- 0x7730
		x"FB",x"F6",x"80",x"01",x"0B",x"00",x"09",x"77", -- 0x7738
		x"E1",x"D1",x"46",x"23",x"5E",x"23",x"CD",x"10", -- 0x7740
		x"75",x"10",x"F9",x"CD",x"21",x"75",x"DA",x"8E", -- 0x7748
		x"74",x"C3",x"A2",x"56",x"40",x"00",x"45",x"14", -- 0x7750
		x"06",x"80",x"11",x"06",x"00",x"FE",x"C7",x"CA", -- 0x7758
		x"AF",x"7A",x"78",x"C3",x"35",x"6C",x"ED",x"5B", -- 0x7760
		x"DC",x"F3",x"D5",x"FE",x"2C",x"28",x"0B",x"CD", -- 0x7768
		x"1C",x"52",x"3C",x"D1",x"57",x"D5",x"2B",x"D7", -- 0x7770
		x"28",x"25",x"CF",x"2C",x"FE",x"2C",x"28",x"0B", -- 0x7778
		x"CD",x"1C",x"52",x"3C",x"D1",x"5F",x"D5",x"2B", -- 0x7780
		x"D7",x"28",x"14",x"CF",x"2C",x"CD",x"1C",x"52", -- 0x7788
		x"A7",x"3E",x"79",x"20",x"01",x"3D",x"F5",x"3E", -- 0x7790
		x"1B",x"DF",x"F1",x"DF",x"3E",x"35",x"DF",x"E3", -- 0x7798
		x"CD",x"C6",x"00",x"E1",x"C9",x"E5",x"21",x"6A", -- 0x77A0
		x"FC",x"18",x"24",x"E5",x"21",x"6D",x"FC",x"18", -- 0x77A8
		x"1E",x"CF",x"45",x"CF",x"52",x"CF",x"FF",x"CF", -- 0x77B0
		x"94",x"E5",x"21",x"7F",x"FC",x"18",x"10",x"3E", -- 0x77B8
		x"04",x"CD",x"08",x"7C",x"2B",x"D7",x"E5",x"16", -- 0x77C0
		x"00",x"21",x"70",x"FC",x"19",x"19",x"19",x"CD", -- 0x77C8
		x"FE",x"77",x"18",x"0E",x"CD",x"1C",x"52",x"3D", -- 0x77D0
		x"FE",x"0A",x"D2",x"5A",x"47",x"7E",x"E5",x"CD", -- 0x77D8
		x"E8",x"77",x"E1",x"F1",x"D7",x"C3",x"12",x"46", -- 0x77E0
		x"16",x"00",x"21",x"CD",x"FB",x"19",x"E5",x"21", -- 0x77E8
		x"49",x"FC",x"19",x"19",x"19",x"CD",x"FE",x"77", -- 0x77F0
		x"7E",x"E6",x"01",x"E1",x"77",x"C9",x"FE",x"95", -- 0x77F8
		x"CA",x"1B",x"63",x"FE",x"EB",x"CA",x"2B",x"63", -- 0x7800
		x"FE",x"90",x"CA",x"31",x"63",x"C3",x"55",x"40", -- 0x7808
		x"CD",x"EA",x"FD",x"01",x"0A",x"00",x"FE",x"CC", -- 0x7810
		x"C8",x"01",x"01",x"0A",x"FE",x"90",x"C8",x"04", -- 0x7818
		x"FE",x"C7",x"C8",x"FE",x"FF",x"D8",x"E5",x"D7", -- 0x7820
		x"FE",x"A3",x"28",x"07",x"FE",x"85",x"28",x"08", -- 0x7828
		x"E1",x"37",x"C9",x"C1",x"01",x"05",x"0C",x"C9", -- 0x7830
		x"D7",x"FE",x"45",x"20",x"F3",x"C1",x"D7",x"CF", -- 0x7838
		x"52",x"CF",x"FF",x"CF",x"94",x"CF",x"EF",x"CD", -- 0x7840
		x"2F",x"54",x"7A",x"B3",x"CA",x"5A",x"47",x"EB", -- 0x7848
		x"22",x"A0",x"FC",x"22",x"A2",x"FC",x"EB",x"01", -- 0x7850
		x"01",x"11",x"2B",x"C9",x"E5",x"47",x"87",x"80", -- 0x7858
		x"6F",x"26",x"00",x"01",x"4D",x"FC",x"09",x"73", -- 0x7860
		x"23",x"72",x"E1",x"C9",x"FE",x"93",x"20",x"3E", -- 0x7868
		x"D7",x"E5",x"21",x"7F",x"F8",x"0E",x"0A",x"06", -- 0x7870
		x"10",x"7E",x"23",x"CD",x"AB",x"00",x"38",x"11", -- 0x7878
		x"05",x"28",x"1B",x"7E",x"23",x"5F",x"CD",x"AB", -- 0x7880
		x"00",x"28",x"06",x"3E",x"01",x"DF",x"7B",x"18", -- 0x7888
		x"0A",x"FE",x"7F",x"28",x"04",x"FE",x"20",x"30", -- 0x7890
		x"02",x"3E",x"20",x"DF",x"10",x"DB",x"CD",x"28", -- 0x7898
		x"73",x"0D",x"20",x"D3",x"E1",x"C9",x"D7",x"C3", -- 0x78A0
		x"CF",x"00",x"D7",x"C3",x"CC",x"00",x"FE",x"28", -- 0x78A8
		x"CA",x"D4",x"77",x"FE",x"95",x"28",x"EF",x"FE", -- 0x78B0
		x"EB",x"28",x"EF",x"CD",x"1C",x"52",x"3D",x"FE", -- 0x78B8
		x"0A",x"D2",x"5A",x"47",x"EB",x"6F",x"26",x"00", -- 0x78C0
		x"29",x"29",x"29",x"29",x"01",x"7F",x"F8",x"09", -- 0x78C8
		x"E5",x"EB",x"CF",x"2C",x"CD",x"64",x"4C",x"E5", -- 0x78D0
		x"CD",x"D0",x"67",x"46",x"23",x"5E",x"23",x"56", -- 0x78D8
		x"E1",x"E3",x"0E",x"0F",x"78",x"A7",x"28",x"0D", -- 0x78E0
		x"1A",x"A7",x"CA",x"5A",x"47",x"77",x"13",x"23", -- 0x78E8
		x"0D",x"28",x"07",x"10",x"F3",x"70",x"23",x"0D", -- 0x78F0
		x"20",x"FB",x"71",x"CD",x"C9",x"00",x"E1",x"C9", -- 0x78F8
		x"D7",x"E5",x"2A",x"9E",x"FC",x"CD",x"36",x"32", -- 0x7900
		x"E1",x"C9",x"D7",x"E5",x"3A",x"DC",x"F3",x"18", -- 0x7908
		x"21",x"CF",x"EF",x"CD",x"2F",x"54",x"ED",x"53", -- 0x7910
		x"9E",x"FC",x"C9",x"D7",x"3E",x"03",x"CD",x"08", -- 0x7918
		x"7C",x"E5",x"3A",x"3F",x"FB",x"1D",x"FA",x"38", -- 0x7920
		x"79",x"0F",x"1D",x"F2",x"29",x"79",x"3E",x"00", -- 0x7928
		x"30",x"01",x"3D",x"CD",x"9A",x"2E",x"E1",x"C9", -- 0x7930
		x"E6",x"07",x"28",x"F7",x"3E",x"FF",x"18",x"F3", -- 0x7938
		x"CD",x"1F",x"52",x"FE",x"03",x"30",x"0A",x"CD", -- 0x7940
		x"D5",x"00",x"18",x"1A",x"CD",x"1F",x"52",x"FE", -- 0x7948
		x"05",x"D2",x"5A",x"47",x"CD",x"D8",x"00",x"C3", -- 0x7950
		x"9A",x"2E",x"CD",x"1F",x"52",x"3D",x"FE",x"0C", -- 0x7958
		x"30",x"EF",x"3C",x"CD",x"DE",x"00",x"C3",x"CF", -- 0x7960
		x"4F",x"CD",x"1F",x"52",x"FE",x"08",x"30",x"E1", -- 0x7968
		x"F5",x"CD",x"DB",x"00",x"47",x"F1",x"E6",x"03", -- 0x7970
		x"3D",x"FE",x"02",x"78",x"38",x"E8",x"18",x"D7", -- 0x7978
		x"01",x"5A",x"47",x"C5",x"ED",x"5B",x"E9",x"F3", -- 0x7980
		x"D5",x"FE",x"2C",x"28",x"0D",x"CD",x"1C",x"52", -- 0x7988
		x"D1",x"FE",x"10",x"D0",x"5F",x"D5",x"2B",x"D7", -- 0x7990
		x"28",x"22",x"CF",x"2C",x"28",x"1E",x"FE",x"2C", -- 0x7998
		x"28",x"0D",x"CD",x"1C",x"52",x"D1",x"FE",x"10", -- 0x79A0
		x"D0",x"57",x"D5",x"2B",x"D7",x"28",x"0D",x"CF", -- 0x79A8
		x"2C",x"CD",x"1C",x"52",x"D1",x"FE",x"10",x"D0", -- 0x79B0
		x"32",x"EB",x"F3",x"D5",x"D1",x"F1",x"E5",x"EB", -- 0x79B8
		x"22",x"E9",x"F3",x"7D",x"32",x"F2",x"F3",x"CD", -- 0x79C0
		x"62",x"00",x"E1",x"C9",x"CD",x"C0",x"FF",x"FE", -- 0x79C8
		x"2C",x"28",x"17",x"CD",x"1C",x"52",x"FE",x"04", -- 0x79D0
		x"D2",x"5A",x"47",x"E5",x"CD",x"5F",x"00",x"3A", -- 0x79D8
		x"B0",x"F3",x"5F",x"CD",x"01",x"52",x"E1",x"2B", -- 0x79E0
		x"D7",x"C8",x"CF",x"2C",x"FE",x"2C",x"28",x"19", -- 0x79E8
		x"CD",x"1C",x"52",x"FE",x"04",x"D2",x"5A",x"47", -- 0x79F0
		x"3A",x"E0",x"F3",x"E6",x"FC",x"B3",x"32",x"E0", -- 0x79F8
		x"F3",x"E5",x"CD",x"69",x"00",x"E1",x"2B",x"D7", -- 0x7A00
		x"C8",x"CF",x"2C",x"FE",x"2C",x"28",x"09",x"CD", -- 0x7A08
		x"1C",x"52",x"32",x"DB",x"F3",x"2B",x"D7",x"C8", -- 0x7A10
		x"CF",x"2C",x"FE",x"2C",x"28",x"06",x"CD",x"2D", -- 0x7A18
		x"7A",x"2B",x"D7",x"C8",x"CF",x"2C",x"CD",x"1C", -- 0x7A20
		x"52",x"32",x"17",x"F4",x"C9",x"CD",x"1C",x"52", -- 0x7A28
		x"3D",x"FE",x"02",x"D2",x"5A",x"47",x"E5",x"01", -- 0x7A30
		x"05",x"00",x"A7",x"21",x"FC",x"F3",x"28",x"01", -- 0x7A38
		x"09",x"11",x"06",x"F4",x"ED",x"B0",x"E1",x"C9", -- 0x7A40
		x"FE",x"24",x"C2",x"AB",x"77",x"3A",x"AF",x"FC", -- 0x7A48
		x"A7",x"CA",x"5A",x"47",x"CD",x"A0",x"7A",x"D5", -- 0x7A50
		x"CD",x"5F",x"4C",x"E3",x"E5",x"CD",x"D0",x"67", -- 0x7A58
		x"23",x"5E",x"23",x"56",x"CD",x"8A",x"00",x"4F", -- 0x7A60
		x"06",x"00",x"2B",x"2B",x"3D",x"BE",x"7E",x"38", -- 0x7A68
		x"0C",x"E1",x"E5",x"F5",x"AF",x"CD",x"56",x"00", -- 0x7A70
		x"F1",x"A7",x"4F",x"06",x"00",x"EB",x"D1",x"C4", -- 0x7A78
		x"5C",x"00",x"E1",x"C9",x"CD",x"9F",x"7A",x"E5", -- 0x7A80
		x"D5",x"CD",x"8A",x"00",x"4F",x"06",x"00",x"C5", -- 0x7A88
		x"CD",x"27",x"66",x"2A",x"99",x"F6",x"EB",x"C1", -- 0x7A90
		x"E1",x"CD",x"59",x"00",x"C3",x"54",x"66",x"D7", -- 0x7A98
		x"CF",x"24",x"3E",x"FF",x"CD",x"08",x"7C",x"E5", -- 0x7AA0
		x"7B",x"CD",x"84",x"00",x"EB",x"E1",x"C9",x"05", -- 0x7AA8
		x"FA",x"5A",x"47",x"3A",x"AF",x"FC",x"A7",x"CA", -- 0x7AB0
		x"5A",x"47",x"D7",x"CD",x"1C",x"52",x"FE",x"20", -- 0x7AB8
		x"D2",x"5A",x"47",x"E5",x"CD",x"87",x"00",x"E3", -- 0x7AC0
		x"CF",x"2C",x"FE",x"2C",x"28",x"2B",x"CD",x"9C", -- 0x7AC8
		x"57",x"E3",x"7B",x"CD",x"4D",x"00",x"78",x"87", -- 0x7AD0
		x"79",x"06",x"00",x"30",x"04",x"C6",x"20",x"06", -- 0x7AD8
		x"80",x"23",x"CD",x"4D",x"00",x"23",x"23",x"CD", -- 0x7AE0
		x"4A",x"00",x"E6",x"0F",x"B0",x"CD",x"4D",x"00", -- 0x7AE8
		x"2B",x"2B",x"2B",x"E3",x"2B",x"D7",x"C1",x"C8", -- 0x7AF0
		x"C5",x"CF",x"2C",x"FE",x"2C",x"28",x"1E",x"CD", -- 0x7AF8
		x"1C",x"52",x"FE",x"10",x"D2",x"5A",x"47",x"E3", -- 0x7B00
		x"23",x"23",x"23",x"CD",x"4A",x"00",x"E6",x"80", -- 0x7B08
		x"B3",x"CD",x"4D",x"00",x"2B",x"2B",x"2B",x"E3", -- 0x7B10
		x"2B",x"D7",x"C1",x"C8",x"C5",x"CF",x"2C",x"CD", -- 0x7B18
		x"1C",x"52",x"CD",x"8A",x"00",x"7B",x"30",x"07", -- 0x7B20
		x"FE",x"40",x"D2",x"5A",x"47",x"87",x"87",x"E3", -- 0x7B28
		x"23",x"23",x"CD",x"4D",x"00",x"E1",x"C9",x"3E", -- 0x7B30
		x"07",x"CD",x"08",x"7C",x"D5",x"CF",x"EF",x"CD", -- 0x7B38
		x"1C",x"52",x"C1",x"47",x"C3",x"47",x"00",x"D7", -- 0x7B40
		x"3E",x"08",x"CD",x"08",x"7C",x"E5",x"16",x"00", -- 0x7B48
		x"21",x"DF",x"F3",x"19",x"7E",x"CD",x"CF",x"4F", -- 0x7B50
		x"E1",x"C9",x"3E",x"13",x"CD",x"08",x"7C",x"16", -- 0x7B58
		x"00",x"D5",x"CF",x"EF",x"CD",x"64",x"4C",x"E3", -- 0x7B60
		x"E5",x"CD",x"FE",x"7B",x"4D",x"44",x"E1",x"7D", -- 0x7B68
		x"F5",x"29",x"EB",x"21",x"A3",x"7B",x"19",x"79", -- 0x7B70
		x"A6",x"20",x"03",x"23",x"78",x"A6",x"C2",x"5A", -- 0x7B78
		x"47",x"21",x"B3",x"F3",x"19",x"71",x"23",x"70", -- 0x7B80
		x"F1",x"1E",x"FF",x"1C",x"D6",x"05",x"30",x"FB", -- 0x7B88
		x"3A",x"AF",x"FC",x"BB",x"CC",x"99",x"7B",x"E1", -- 0x7B90
		x"C9",x"3D",x"FA",x"78",x"00",x"CA",x"7E",x"00", -- 0x7B98
		x"C3",x"81",x"00",x"FF",x"03",x"3F",x"00",x"FF", -- 0x7BA0
		x"07",x"7F",x"00",x"FF",x"07",x"FF",x"03",x"3F", -- 0x7BA8
		x"00",x"FF",x"07",x"7F",x"00",x"FF",x"07",x"FF", -- 0x7BB0
		x"03",x"FF",x"1F",x"FF",x"1F",x"7F",x"00",x"FF", -- 0x7BB8
		x"07",x"FF",x"03",x"3F",x"00",x"FF",x"07",x"7F", -- 0x7BC0
		x"00",x"FF",x"07",x"D7",x"3E",x"13",x"CD",x"08", -- 0x7BC8
		x"7C",x"E5",x"16",x"00",x"21",x"B3",x"F3",x"19", -- 0x7BD0
		x"19",x"7E",x"23",x"66",x"6F",x"CD",x"36",x"32", -- 0x7BD8
		x"E1",x"C9",x"CD",x"64",x"4C",x"E5",x"CD",x"FE", -- 0x7BE0
		x"7B",x"E3",x"CF",x"2C",x"CD",x"1C",x"52",x"E3", -- 0x7BE8
		x"CD",x"4D",x"00",x"E1",x"C9",x"CD",x"FE",x"7B", -- 0x7BF0
		x"CD",x"4A",x"00",x"C3",x"CF",x"4F",x"CD",x"8A", -- 0x7BF8
		x"2F",x"11",x"00",x"40",x"E7",x"D8",x"18",x"6B", -- 0x7C00
		x"F5",x"CF",x"28",x"CD",x"1C",x"52",x"F1",x"BB", -- 0x7C08
		x"38",x"61",x"CF",x"29",x"7B",x"C9",x"CD",x"EF", -- 0x7C10
		x"FD",x"18",x"58",x"CD",x"F4",x"FD",x"18",x"53", -- 0x7C18
		x"CD",x"F9",x"FD",x"18",x"4E",x"CD",x"FE",x"FD", -- 0x7C20
		x"18",x"49",x"CD",x"03",x"FE",x"18",x"44",x"CD", -- 0x7C28
		x"08",x"FE",x"18",x"3F",x"CD",x"0D",x"FE",x"18", -- 0x7C30
		x"3A",x"CD",x"12",x"FE",x"18",x"35",x"CD",x"17", -- 0x7C38
		x"FE",x"18",x"30",x"CD",x"1C",x"FE",x"18",x"2B", -- 0x7C40
		x"CD",x"21",x"FE",x"18",x"26",x"CD",x"26",x"FE", -- 0x7C48
		x"18",x"21",x"CD",x"2B",x"FE",x"18",x"1C",x"CD", -- 0x7C50
		x"30",x"FE",x"18",x"17",x"CD",x"35",x"FE",x"18", -- 0x7C58
		x"12",x"CD",x"3A",x"FE",x"18",x"0D",x"CD",x"3F", -- 0x7C60
		x"FE",x"18",x"08",x"CD",x"44",x"FE",x"18",x"03", -- 0x7C68
		x"CD",x"49",x"FE",x"C3",x"5A",x"47",x"31",x"76", -- 0x7C70
		x"F3",x"01",x"2F",x"02",x"11",x"9B",x"FD",x"21", -- 0x7C78
		x"9A",x"FD",x"36",x"C9",x"ED",x"B0",x"21",x"80", -- 0x7C80
		x"F3",x"22",x"4A",x"FC",x"CD",x"5D",x"7D",x"22", -- 0x7C88
		x"48",x"FC",x"01",x"90",x"00",x"11",x"80",x"F3", -- 0x7C90
		x"21",x"27",x"7F",x"ED",x"B0",x"CD",x"3E",x"00", -- 0x7C98
		x"AF",x"32",x"60",x"F6",x"32",x"7C",x"F8",x"3E", -- 0x7CA0
		x"2C",x"32",x"5D",x"F5",x"3E",x"3A",x"32",x"1E", -- 0x7CA8
		x"F4",x"2A",x"04",x"00",x"22",x"20",x"F9",x"21", -- 0x7CB0
		x"E4",x"F6",x"22",x"4C",x"F7",x"22",x"74",x"F6", -- 0x7CB8
		x"01",x"C8",x"00",x"09",x"22",x"72",x"F6",x"3E", -- 0x7CC0
		x"01",x"32",x"C3",x"F6",x"CD",x"6B",x"7E",x"CD", -- 0x7CC8
		x"E5",x"62",x"2A",x"48",x"FC",x"AF",x"77",x"23", -- 0x7CD0
		x"22",x"76",x"F6",x"CD",x"87",x"62",x"CD",x"3B", -- 0x7CD8
		x"00",x"CD",x"6F",x"00",x"CD",x"69",x"00",x"21", -- 0x7CE0
		x"0B",x"0A",x"22",x"DC",x"F3",x"21",x"D8",x"7E", -- 0x7CE8
		x"CD",x"78",x"66",x"21",x"0C",x"0A",x"22",x"DC", -- 0x7CF0
		x"F3",x"21",x"E4",x"7E",x"CD",x"78",x"66",x"21", -- 0x7CF8
		x"0E",x"02",x"22",x"DC",x"F3",x"21",x"FD",x"7E", -- 0x7D00
		x"CD",x"78",x"66",x"06",x"06",x"2B",x"7D",x"B4", -- 0x7D08
		x"20",x"FB",x"10",x"F9",x"CD",x"75",x"7D",x"2A", -- 0x7D10
		x"48",x"FC",x"AF",x"77",x"23",x"22",x"76",x"F6", -- 0x7D18
		x"CD",x"87",x"62",x"CD",x"29",x"7D",x"C3",x"1F", -- 0x7D20
		x"41",x"3E",x"FF",x"32",x"DE",x"F3",x"CD",x"6C", -- 0x7D28
		x"00",x"21",x"F2",x"7E",x"CD",x"78",x"66",x"21", -- 0x7D30
		x"E4",x"7E",x"CD",x"78",x"66",x"21",x"FD",x"7E", -- 0x7D38
		x"CD",x"78",x"66",x"2A",x"C2",x"F6",x"EB",x"2A", -- 0x7D40
		x"74",x"F6",x"7D",x"93",x"6F",x"7C",x"9A",x"67", -- 0x7D48
		x"01",x"F2",x"FF",x"09",x"CD",x"12",x"34",x"21", -- 0x7D50
		x"1B",x"7F",x"C3",x"78",x"66",x"21",x"00",x"EF", -- 0x7D58
		x"7E",x"2F",x"77",x"BE",x"2F",x"77",x"20",x"09", -- 0x7D60
		x"2C",x"20",x"F5",x"7C",x"3D",x"F0",x"67",x"18", -- 0x7D68
		x"EF",x"2E",x"00",x"24",x"C9",x"F3",x"0E",x"00", -- 0x7D70
		x"11",x"C1",x"FC",x"21",x"C9",x"FC",x"1A",x"B1", -- 0x7D78
		x"4F",x"D5",x"23",x"E5",x"21",x"00",x"40",x"CD", -- 0x7D80
		x"1A",x"7E",x"E5",x"21",x"41",x"42",x"E7",x"E1", -- 0x7D88
		x"06",x"00",x"20",x"2A",x"CD",x"1A",x"7E",x"E5", -- 0x7D90
		x"C5",x"D5",x"DD",x"E1",x"79",x"F5",x"FD",x"E1", -- 0x7D98
		x"C4",x"1C",x"00",x"C1",x"E1",x"CD",x"1A",x"7E", -- 0x7DA0
		x"C6",x"FF",x"CB",x"18",x"CD",x"1A",x"7E",x"C6", -- 0x7DA8
		x"FF",x"CB",x"18",x"CD",x"1A",x"7E",x"C6",x"FF", -- 0x7DB0
		x"CB",x"18",x"11",x"F8",x"FF",x"19",x"E3",x"70", -- 0x7DB8
		x"23",x"E3",x"11",x"FE",x"3F",x"19",x"7C",x"FE", -- 0x7DC0
		x"C0",x"38",x"BC",x"E1",x"23",x"79",x"A7",x"11", -- 0x7DC8
		x"0C",x"00",x"F2",x"E0",x"7D",x"C6",x"04",x"4F", -- 0x7DD0
		x"FE",x"90",x"38",x"A6",x"E6",x"03",x"4F",x"3E", -- 0x7DD8
		x"19",x"D1",x"13",x"0C",x"79",x"FE",x"04",x"38", -- 0x7DE0
		x"95",x"21",x"C9",x"FC",x"06",x"40",x"7E",x"87", -- 0x7DE8
		x"38",x"04",x"23",x"10",x"F9",x"C9",x"CD",x"2A", -- 0x7DF0
		x"7E",x"CD",x"24",x"00",x"2A",x"C2",x"F6",x"11", -- 0x7DF8
		x"00",x"C0",x"E7",x"30",x"04",x"EB",x"22",x"C2", -- 0x7E00
		x"F6",x"2A",x"08",x"80",x"23",x"22",x"76",x"F6", -- 0x7E08
		x"7C",x"32",x"B1",x"FB",x"CD",x"9A",x"62",x"C3", -- 0x7E10
		x"01",x"46",x"CD",x"1E",x"7E",x"5A",x"79",x"C5", -- 0x7E18
		x"D5",x"CD",x"0C",x"00",x"D1",x"C1",x"57",x"B3", -- 0x7E20
		x"23",x"C9",x"3E",x"40",x"90",x"47",x"26",x"00", -- 0x7E28
		x"1F",x"CB",x"1C",x"1F",x"CB",x"1C",x"1F",x"1F", -- 0x7E30
		x"E6",x"03",x"4F",x"78",x"06",x"00",x"E5",x"21", -- 0x7E38
		x"C1",x"FC",x"09",x"E6",x"0C",x"B1",x"4F",x"7E", -- 0x7E40
		x"E1",x"B1",x"C9",x"CF",x"B7",x"CF",x"EF",x"CD", -- 0x7E48
		x"1C",x"52",x"C2",x"55",x"40",x"FE",x"10",x"D2", -- 0x7E50
		x"5A",x"47",x"22",x"A7",x"F6",x"F5",x"CD",x"1C", -- 0x7E58
		x"6C",x"F1",x"CD",x"6B",x"7E",x"CD",x"A7",x"62", -- 0x7E60
		x"C3",x"01",x"46",x"F5",x"2A",x"4A",x"FC",x"11", -- 0x7E68
		x"F5",x"FE",x"19",x"3D",x"F2",x"72",x"7E",x"EB", -- 0x7E70
		x"2A",x"74",x"F6",x"44",x"4D",x"2A",x"72",x"F6", -- 0x7E78
		x"7D",x"91",x"6F",x"7C",x"98",x"67",x"F1",x"E5", -- 0x7E80
		x"F5",x"01",x"8C",x"00",x"09",x"44",x"4D",x"2A", -- 0x7E88
		x"C2",x"F6",x"09",x"E7",x"D2",x"75",x"62",x"F1", -- 0x7E90
		x"32",x"5F",x"F8",x"6B",x"62",x"22",x"60",x"F8", -- 0x7E98
		x"2B",x"2B",x"22",x"72",x"F6",x"C1",x"7D",x"91", -- 0x7EA0
		x"6F",x"7C",x"98",x"67",x"22",x"74",x"F6",x"2B", -- 0x7EA8
		x"2B",x"C1",x"F9",x"C5",x"3A",x"5F",x"F8",x"6F", -- 0x7EB0
		x"2C",x"26",x"00",x"29",x"19",x"EB",x"D5",x"01", -- 0x7EB8
		x"09",x"01",x"73",x"23",x"72",x"23",x"EB",x"36", -- 0x7EC0
		x"00",x"09",x"EB",x"3D",x"F2",x"C2",x"7E",x"E1", -- 0x7EC8
		x"01",x"09",x"00",x"09",x"22",x"62",x"F8",x"C9", -- 0x7ED0
		x"4D",x"53",x"58",x"20",x"20",x"73",x"79",x"73", -- 0x7ED8
		x"74",x"65",x"6D",x"00",x"76",x"65",x"72",x"73", -- 0x7EE0
		x"69",x"6F",x"6E",x"20",x"31",x"2E",x"30",x"0D", -- 0x7EE8
		x"0A",x"00",x"4D",x"53",x"58",x"20",x"42",x"41", -- 0x7EF0
		x"53",x"49",x"43",x"20",x"00",x"43",x"6F",x"70", -- 0x7EF8
		x"79",x"72",x"69",x"67",x"68",x"74",x"20",x"31", -- 0x7F00
		x"39",x"38",x"33",x"20",x"62",x"79",x"20",x"4D", -- 0x7F08
		x"69",x"63",x"72",x"6F",x"73",x"6F",x"66",x"74", -- 0x7F10
		x"0D",x"0A",x"00",x"20",x"42",x"79",x"74",x"65", -- 0x7F18
		x"73",x"20",x"66",x"72",x"65",x"65",x"00",x"D3", -- 0x7F20
		x"A8",x"5E",x"18",x"03",x"D3",x"A8",x"73",x"7A", -- 0x7F28
		x"D3",x"A8",x"C9",x"D3",x"A8",x"08",x"CD",x"98", -- 0x7F30
		x"F3",x"08",x"F1",x"D3",x"A8",x"08",x"C9",x"DD", -- 0x7F38
		x"E9",x"5A",x"47",x"5A",x"47",x"5A",x"47",x"5A", -- 0x7F40
		x"47",x"5A",x"47",x"5A",x"47",x"5A",x"47",x"5A", -- 0x7F48
		x"47",x"5A",x"47",x"5A",x"47",x"25",x"1D",x"1D", -- 0x7F50
		x"18",x"0E",x"00",x"00",x"00",x"00",x"00",x"08", -- 0x7F58
		x"00",x"00",x"00",x"00",x"00",x"18",x"00",x"20", -- 0x7F60
		x"00",x"00",x"00",x"1B",x"00",x"38",x"00",x"18", -- 0x7F68
		x"00",x"20",x"00",x"00",x"00",x"1B",x"00",x"38", -- 0x7F70
		x"00",x"08",x"00",x"00",x"00",x"00",x"00",x"1B", -- 0x7F78
		x"00",x"38",x"01",x"01",x"01",x"00",x"00",x"E0", -- 0x7F80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF", -- 0x7F88
		x"0F",x"04",x"04",x"C3",x"00",x"00",x"C3",x"00", -- 0x7F90
		x"00",x"0F",x"59",x"F9",x"FF",x"01",x"32",x"F0", -- 0x7F98
		x"FB",x"F0",x"FB",x"53",x"5C",x"26",x"2D",x"0F", -- 0x7FA0
		x"25",x"2D",x"0E",x"16",x"1F",x"53",x"5C",x"26", -- 0x7FA8
		x"2D",x"0F",x"00",x"01",x"00",x"01",x"3A",x"11", -- 0x7FB0
		x"89",x"FD",x"A7",x"C0",x"04",x"C9",x"CD",x"CB", -- 0x7FB8
		x"7F",x"5E",x"18",x"04",x"CD",x"CB",x"7F",x"73", -- 0x7FC0
		x"78",x"18",x"0E",x"0F",x"0F",x"E6",x"03",x"57", -- 0x7FC8
		x"3A",x"FF",x"FF",x"2F",x"47",x"E6",x"FC",x"B2", -- 0x7FD0
		x"57",x"32",x"FF",x"FF",x"7B",x"C9",x"00",x"00", -- 0x7FD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7FE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7FE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x7FF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"  -- 0x7FF8
	);

begin

	process(clk)
	begin
		if rising_edge(clk) then
			data <= ROM(to_integer(unsigned(addr)));
		end if;
	end process;
end RTL;
