-- generated with romgen v3.0 by MikeJ
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity ipl_rom is
	port (
		clk		: in    std_logic;
		addr		: in    std_logic_vector(12 downto 0);
		data		: out   std_logic_vector(7 downto 0)
	);
end;

architecture rtl of ipl_rom is

	type ROM_ARRAY is array(0 to 8191) of std_logic_vector(7 downto 0);
	constant ROM : ROM_ARRAY := (
		x"F3",x"ED",x"56",x"C3",x"80",x"00",x"FF",x"FF", -- 0x0000
		x"ED",x"4D",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0008
		x"ED",x"4D",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0010
		x"ED",x"4D",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0018
		x"ED",x"4D",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0020
		x"ED",x"4D",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0028
		x"ED",x"4D",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0030
		x"ED",x"4D",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0038
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0040
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0048
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0050
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0058
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"ED",x"45", -- 0x0060
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0068
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0070
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0078
		x"31",x"FF",x"7F",x"CD",x"7A",x"1B",x"CD",x"75", -- 0x0080
		x"01",x"C3",x"00",x"01",x"FF",x"FF",x"FF",x"FF", -- 0x0088
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0090
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0098
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00A8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00F8
		x"76",x"18",x"FD",x"21",x"03",x"00",x"39",x"4E", -- 0x0100
		x"23",x"46",x"C5",x"CD",x"C1",x"19",x"F1",x"CB", -- 0x0108
		x"3C",x"CB",x"1D",x"55",x"3E",x"10",x"92",x"57", -- 0x0110
		x"21",x"02",x"00",x"39",x"7E",x"F5",x"33",x"D5", -- 0x0118
		x"33",x"CD",x"C5",x"18",x"F1",x"21",x"03",x"00", -- 0x0120
		x"39",x"4E",x"23",x"46",x"C5",x"CD",x"AE",x"19", -- 0x0128
		x"F1",x"C9",x"28",x"20",x"20",x"20",x"20",x"20", -- 0x0130
		x"20",x"20",x"20",x"4D",x"53",x"58",x"31",x"20", -- 0x0138
		x"46",x"50",x"47",x"41",x"20",x"4C",x"4F",x"41", -- 0x0140
		x"44",x"45",x"52",x"20",x"20",x"20",x"20",x"20", -- 0x0148
		x"20",x"20",x"20",x"00",x"3E",x"FF",x"D3",x"9E", -- 0x0150
		x"21",x"01",x"0F",x"E5",x"3E",x"06",x"F5",x"33", -- 0x0158
		x"CD",x"4B",x"18",x"F1",x"33",x"C1",x"E1",x"E5", -- 0x0160
		x"C5",x"E5",x"3E",x"0C",x"F5",x"33",x"CD",x"03", -- 0x0168
		x"01",x"F1",x"33",x"18",x"FE",x"21",x"CB",x"FD", -- 0x0170
		x"39",x"F9",x"21",x"33",x"02",x"39",x"AF",x"77", -- 0x0178
		x"23",x"77",x"CD",x"BD",x"17",x"21",x"01",x"0F", -- 0x0180
		x"E5",x"3E",x"04",x"F5",x"33",x"CD",x"4B",x"18", -- 0x0188
		x"33",x"21",x"33",x"01",x"E3",x"CD",x"AE",x"19", -- 0x0190
		x"F1",x"3A",x"32",x"01",x"D3",x"40",x"3E",x"12", -- 0x0198
		x"D3",x"48",x"3E",x"01",x"D3",x"49",x"3E",x"00", -- 0x01A0
		x"D3",x"48",x"DB",x"49",x"4F",x"3E",x"01",x"D3", -- 0x01A8
		x"48",x"21",x"00",x"00",x"39",x"FD",x"21",x"2F", -- 0x01B0
		x"02",x"FD",x"39",x"FD",x"75",x"00",x"FD",x"74", -- 0x01B8
		x"01",x"06",x"00",x"FD",x"21",x"2F",x"02",x"FD", -- 0x01C0
		x"39",x"FD",x"7E",x"00",x"80",x"5F",x"FD",x"7E", -- 0x01C8
		x"01",x"CE",x"00",x"57",x"DB",x"49",x"12",x"1A", -- 0x01D0
		x"B7",x"28",x"06",x"04",x"78",x"D6",x"14",x"38", -- 0x01D8
		x"E2",x"3E",x"02",x"D3",x"48",x"DB",x"49",x"47", -- 0x01E0
		x"C5",x"21",x"00",x"03",x"E5",x"CD",x"C5",x"18", -- 0x01E8
		x"F1",x"C1",x"21",x"13",x"08",x"C5",x"E5",x"CD", -- 0x01F0
		x"AE",x"19",x"F1",x"C1",x"79",x"C6",x"30",x"C5", -- 0x01F8
		x"F5",x"33",x"CD",x"3B",x"19",x"33",x"C1",x"21", -- 0x0200
		x"1C",x"08",x"C5",x"E5",x"CD",x"AE",x"19",x"F1", -- 0x0208
		x"C1",x"21",x"2F",x"02",x"39",x"7E",x"23",x"66", -- 0x0210
		x"6F",x"C5",x"E5",x"CD",x"AE",x"19",x"F1",x"C1", -- 0x0218
		x"21",x"20",x"08",x"C5",x"E5",x"CD",x"AE",x"19", -- 0x0220
		x"F1",x"C1",x"78",x"07",x"07",x"07",x"07",x"E6", -- 0x0228
		x"0F",x"C6",x"30",x"C5",x"F5",x"33",x"CD",x"3B", -- 0x0230
		x"19",x"33",x"3E",x"2E",x"F5",x"33",x"CD",x"3B", -- 0x0238
		x"19",x"33",x"C1",x"78",x"E6",x"0F",x"C6",x"30", -- 0x0240
		x"C5",x"F5",x"33",x"CD",x"3B",x"19",x"33",x"C1", -- 0x0248
		x"21",x"2B",x"08",x"C5",x"E5",x"CD",x"AE",x"19", -- 0x0250
		x"F1",x"C1",x"21",x"2E",x"08",x"C5",x"E5",x"CD", -- 0x0258
		x"AE",x"19",x"F1",x"CD",x"BE",x"0A",x"7D",x"C1", -- 0x0260
		x"B7",x"20",x"0A",x"21",x"45",x"08",x"C5",x"E5", -- 0x0268
		x"CD",x"54",x"01",x"F1",x"C1",x"C5",x"CD",x"17", -- 0x0270
		x"0F",x"C1",x"7C",x"B5",x"20",x"0A",x"21",x"66", -- 0x0278
		x"08",x"C5",x"E5",x"CD",x"54",x"01",x"F1",x"C1", -- 0x0280
		x"21",x"78",x"08",x"C5",x"E5",x"CD",x"AE",x"19", -- 0x0288
		x"F1",x"2A",x"28",x"44",x"E5",x"CD",x"A6",x"13", -- 0x0290
		x"F1",x"C1",x"7C",x"B5",x"20",x"0A",x"21",x"92", -- 0x0298
		x"08",x"C5",x"E5",x"CD",x"54",x"01",x"F1",x"C1", -- 0x02A0
		x"21",x"15",x"02",x"39",x"FD",x"21",x"2F",x"02", -- 0x02A8
		x"FD",x"39",x"FD",x"75",x"00",x"FD",x"74",x"01", -- 0x02B0
		x"FD",x"5E",x"00",x"FD",x"56",x"01",x"C5",x"2A", -- 0x02B8
		x"2A",x"44",x"E5",x"D5",x"CD",x"3C",x"12",x"F1", -- 0x02C0
		x"F1",x"C1",x"7C",x"B5",x"20",x"0A",x"21",x"B2", -- 0x02C8
		x"08",x"C5",x"E5",x"CD",x"54",x"01",x"F1",x"C1", -- 0x02D0
		x"21",x"31",x"02",x"39",x"FD",x"21",x"2F",x"02", -- 0x02D8
		x"FD",x"39",x"FD",x"7E",x"00",x"C6",x"01",x"77", -- 0x02E0
		x"FD",x"7E",x"01",x"CE",x"00",x"23",x"77",x"21", -- 0x02E8
		x"31",x"02",x"39",x"7E",x"23",x"66",x"6F",x"56", -- 0x02F0
		x"23",x"5E",x"23",x"46",x"23",x"66",x"7A",x"D6", -- 0x02F8
		x"03",x"7B",x"DE",x"00",x"78",x"DE",x"00",x"7C", -- 0x0300
		x"DE",x"00",x"30",x"0A",x"21",x"C9",x"08",x"C5", -- 0x0308
		x"E5",x"CD",x"54",x"01",x"F1",x"C1",x"21",x"15", -- 0x0310
		x"00",x"39",x"FD",x"21",x"2D",x"02",x"FD",x"39", -- 0x0318
		x"FD",x"75",x"00",x"FD",x"74",x"01",x"FD",x"5E", -- 0x0320
		x"00",x"FD",x"56",x"01",x"21",x"2F",x"02",x"39", -- 0x0328
		x"7E",x"23",x"66",x"6F",x"C5",x"D5",x"E5",x"CD", -- 0x0330
		x"99",x"12",x"F1",x"F1",x"C1",x"7C",x"B5",x"20", -- 0x0338
		x"0A",x"21",x"DC",x"08",x"C5",x"E5",x"CD",x"54", -- 0x0340
		x"01",x"F1",x"C1",x"21",x"2D",x"02",x"39",x"7E", -- 0x0348
		x"23",x"66",x"6F",x"7E",x"D6",x"31",x"20",x"04", -- 0x0350
		x"1E",x"01",x"18",x"02",x"1E",x"00",x"21",x"2D", -- 0x0358
		x"02",x"39",x"7E",x"23",x"66",x"6F",x"23",x"7E", -- 0x0360
		x"D6",x"31",x"20",x"04",x"16",x"02",x"18",x"02", -- 0x0368
		x"16",x"00",x"21",x"2D",x"02",x"39",x"7E",x"23", -- 0x0370
		x"66",x"6F",x"23",x"23",x"7E",x"FD",x"21",x"22", -- 0x0378
		x"02",x"FD",x"39",x"FD",x"77",x"00",x"FD",x"7E", -- 0x0380
		x"00",x"D6",x"45",x"28",x"21",x"FD",x"7E",x"00", -- 0x0388
		x"D6",x"42",x"28",x"1A",x"FD",x"7E",x"00",x"D6", -- 0x0390
		x"46",x"28",x"13",x"FD",x"7E",x"00",x"D6",x"53", -- 0x0398
		x"28",x"0C",x"21",x"F7",x"08",x"C5",x"D5",x"E5", -- 0x03A0
		x"CD",x"54",x"01",x"F1",x"D1",x"C1",x"21",x"2D", -- 0x03A8
		x"02",x"39",x"7E",x"23",x"66",x"6F",x"23",x"23", -- 0x03B0
		x"23",x"7E",x"D6",x"50",x"20",x"04",x"06",x"02", -- 0x03B8
		x"18",x"02",x"06",x"00",x"21",x"2D",x"02",x"39", -- 0x03C0
		x"7E",x"23",x"66",x"6F",x"23",x"23",x"23",x"23", -- 0x03C8
		x"7E",x"D6",x"31",x"20",x"04",x"3E",x"01",x"18", -- 0x03D0
		x"02",x"3E",x"00",x"FD",x"21",x"28",x"02",x"FD", -- 0x03D8
		x"39",x"FD",x"77",x"00",x"78",x"D3",x"99",x"3E", -- 0x03E0
		x"89",x"D3",x"99",x"3E",x"10",x"D3",x"48",x"7A", -- 0x03E8
		x"B3",x"D3",x"49",x"21",x"07",x"09",x"C5",x"D5", -- 0x03F0
		x"E5",x"CD",x"AE",x"19",x"F1",x"D1",x"C1",x"16", -- 0x03F8
		x"00",x"7A",x"D6",x"0F",x"28",x"18",x"21",x"FF", -- 0x0400
		x"3F",x"72",x"E5",x"D5",x"C5",x"21",x"00",x"80", -- 0x0408
		x"11",x"01",x"80",x"01",x"FF",x"3F",x"3E",x"00", -- 0x0410
		x"77",x"ED",x"B0",x"C1",x"D1",x"E1",x"14",x"7A", -- 0x0418
		x"D6",x"20",x"38",x"DD",x"21",x"19",x"09",x"C5", -- 0x0420
		x"D5",x"E5",x"CD",x"AE",x"19",x"F1",x"D1",x"C1", -- 0x0428
		x"79",x"FE",x"05",x"28",x"05",x"D6",x"06",x"C2", -- 0x0430
		x"10",x"05",x"21",x"1E",x"09",x"D5",x"E5",x"CD", -- 0x0438
		x"AE",x"19",x"F1",x"D1",x"21",x"2F",x"02",x"39", -- 0x0440
		x"4E",x"23",x"46",x"D5",x"2A",x"2E",x"44",x"E5", -- 0x0448
		x"C5",x"CD",x"3C",x"12",x"F1",x"F1",x"4D",x"D1", -- 0x0450
		x"7C",x"B1",x"20",x"0A",x"21",x"35",x"09",x"D5", -- 0x0458
		x"E5",x"CD",x"54",x"01",x"F1",x"D1",x"21",x"31", -- 0x0460
		x"02",x"39",x"7E",x"23",x"66",x"6F",x"56",x"23", -- 0x0468
		x"46",x"23",x"4E",x"23",x"66",x"7A",x"B7",x"20", -- 0x0470
		x"0B",x"78",x"D6",x"80",x"20",x"06",x"B1",x"20", -- 0x0478
		x"03",x"B4",x"28",x"0A",x"21",x"4E",x"09",x"D5", -- 0x0480
		x"E5",x"CD",x"54",x"01",x"F1",x"D1",x"21",x"2F", -- 0x0488
		x"02",x"39",x"7E",x"FD",x"21",x"2B",x"02",x"FD", -- 0x0490
		x"39",x"FD",x"77",x"00",x"21",x"30",x"02",x"39", -- 0x0498
		x"7E",x"FD",x"21",x"2B",x"02",x"FD",x"39",x"FD", -- 0x04A0
		x"77",x"01",x"16",x"1E",x"21",x"FF",x"3F",x"72", -- 0x04A8
		x"01",x"00",x"80",x"FD",x"21",x"14",x"00",x"FD", -- 0x04B0
		x"39",x"FD",x"36",x"00",x"00",x"21",x"2B",x"02", -- 0x04B8
		x"39",x"7E",x"23",x"66",x"6F",x"C5",x"D5",x"C5", -- 0x04C0
		x"E5",x"CD",x"99",x"12",x"F1",x"F1",x"D1",x"C1", -- 0x04C8
		x"7C",x"B5",x"20",x"0C",x"21",x"6F",x"09",x"C5", -- 0x04D0
		x"D5",x"E5",x"CD",x"54",x"01",x"F1",x"D1",x"C1", -- 0x04D8
		x"21",x"00",x"02",x"09",x"4D",x"44",x"FD",x"21", -- 0x04E0
		x"14",x"00",x"FD",x"39",x"FD",x"34",x"00",x"FD", -- 0x04E8
		x"7E",x"00",x"D6",x"20",x"38",x"C7",x"D5",x"3E", -- 0x04F0
		x"2E",x"F5",x"33",x"CD",x"3B",x"19",x"33",x"D1", -- 0x04F8
		x"14",x"7A",x"D6",x"20",x"38",x"A6",x"21",x"19", -- 0x0500
		x"09",x"D5",x"E5",x"CD",x"AE",x"19",x"F1",x"D1", -- 0x0508
		x"1D",x"C2",x"1C",x"06",x"21",x"88",x"09",x"E5", -- 0x0510
		x"CD",x"AE",x"19",x"F1",x"21",x"2F",x"02",x"39", -- 0x0518
		x"5E",x"23",x"56",x"2A",x"2C",x"44",x"E5",x"D5", -- 0x0520
		x"CD",x"3C",x"12",x"F1",x"F1",x"4D",x"7C",x"B1", -- 0x0528
		x"20",x"08",x"21",x"9D",x"09",x"E5",x"CD",x"54", -- 0x0530
		x"01",x"F1",x"21",x"31",x"02",x"39",x"7E",x"23", -- 0x0538
		x"66",x"6F",x"56",x"23",x"5E",x"23",x"46",x"23", -- 0x0540
		x"66",x"7A",x"B7",x"20",x"0B",x"B3",x"20",x"08", -- 0x0548
		x"78",x"D6",x"02",x"20",x"03",x"B4",x"28",x"08", -- 0x0550
		x"21",x"B4",x"09",x"E5",x"CD",x"54",x"01",x"F1", -- 0x0558
		x"21",x"2F",x"02",x"39",x"7E",x"FD",x"21",x"2B", -- 0x0560
		x"02",x"FD",x"39",x"FD",x"77",x"00",x"21",x"30", -- 0x0568
		x"02",x"39",x"7E",x"FD",x"21",x"2B",x"02",x"FD", -- 0x0570
		x"39",x"FD",x"77",x"01",x"FD",x"21",x"27",x"02", -- 0x0578
		x"FD",x"39",x"FD",x"36",x"00",x"00",x"21",x"FF", -- 0x0580
		x"3F",x"FD",x"21",x"27",x"02",x"FD",x"39",x"FD", -- 0x0588
		x"7E",x"00",x"77",x"21",x"23",x"02",x"39",x"36", -- 0x0590
		x"00",x"23",x"36",x"80",x"FD",x"21",x"14",x"00", -- 0x0598
		x"FD",x"39",x"FD",x"36",x"00",x"00",x"21",x"2B", -- 0x05A0
		x"02",x"39",x"7E",x"23",x"66",x"6F",x"FD",x"21", -- 0x05A8
		x"23",x"02",x"FD",x"39",x"FD",x"4E",x"00",x"FD", -- 0x05B0
		x"46",x"01",x"C5",x"E5",x"CD",x"99",x"12",x"F1", -- 0x05B8
		x"F1",x"FD",x"21",x"29",x"02",x"FD",x"39",x"FD", -- 0x05C0
		x"74",x"01",x"FD",x"75",x"00",x"21",x"2A",x"02", -- 0x05C8
		x"39",x"7E",x"2B",x"B6",x"20",x"08",x"21",x"D5", -- 0x05D0
		x"09",x"E5",x"CD",x"54",x"01",x"F1",x"21",x"23", -- 0x05D8
		x"02",x"39",x"7E",x"C6",x"00",x"77",x"23",x"7E", -- 0x05E0
		x"CE",x"02",x"77",x"FD",x"21",x"14",x"00",x"FD", -- 0x05E8
		x"39",x"FD",x"34",x"00",x"FD",x"7E",x"00",x"D6", -- 0x05F0
		x"20",x"38",x"AB",x"3E",x"2E",x"F5",x"33",x"CD", -- 0x05F8
		x"3B",x"19",x"33",x"FD",x"21",x"27",x"02",x"FD", -- 0x0600
		x"39",x"FD",x"34",x"00",x"FD",x"7E",x"00",x"D6", -- 0x0608
		x"08",x"DA",x"86",x"05",x"21",x"19",x"09",x"E5", -- 0x0610
		x"CD",x"AE",x"19",x"F1",x"FD",x"21",x"22",x"02", -- 0x0618
		x"FD",x"39",x"FD",x"7E",x"00",x"FE",x"42",x"28", -- 0x0620
		x"22",x"FE",x"45",x"28",x"0A",x"FE",x"46",x"28", -- 0x0628
		x"2E",x"D6",x"53",x"28",x"3E",x"18",x"4E",x"21", -- 0x0630
		x"30",x"44",x"7E",x"FD",x"21",x"33",x"02",x"FD", -- 0x0638
		x"39",x"FD",x"77",x"00",x"23",x"7E",x"FD",x"77", -- 0x0640
		x"01",x"18",x"3A",x"21",x"32",x"44",x"7E",x"FD", -- 0x0648
		x"21",x"33",x"02",x"FD",x"39",x"FD",x"77",x"00", -- 0x0650
		x"23",x"7E",x"FD",x"77",x"01",x"18",x"26",x"21", -- 0x0658
		x"34",x"44",x"7E",x"FD",x"21",x"33",x"02",x"FD", -- 0x0660
		x"39",x"FD",x"77",x"00",x"23",x"7E",x"FD",x"77", -- 0x0668
		x"01",x"18",x"12",x"21",x"36",x"44",x"7E",x"FD", -- 0x0670
		x"21",x"33",x"02",x"FD",x"39",x"FD",x"77",x"00", -- 0x0678
		x"23",x"7E",x"FD",x"77",x"01",x"21",x"F0",x"09", -- 0x0680
		x"E5",x"CD",x"AE",x"19",x"F1",x"21",x"2F",x"02", -- 0x0688
		x"39",x"7E",x"23",x"66",x"6F",x"FD",x"21",x"33", -- 0x0690
		x"02",x"FD",x"39",x"FD",x"4E",x"00",x"FD",x"46", -- 0x0698
		x"01",x"C5",x"E5",x"CD",x"3C",x"12",x"F1",x"F1", -- 0x06A0
		x"7C",x"B5",x"20",x"08",x"21",x"01",x"0A",x"E5", -- 0x06A8
		x"CD",x"54",x"01",x"F1",x"21",x"31",x"02",x"39", -- 0x06B0
		x"7E",x"23",x"66",x"6F",x"56",x"23",x"5E",x"23", -- 0x06B8
		x"46",x"23",x"6E",x"7A",x"B7",x"20",x"0B",x"7B", -- 0x06C0
		x"D6",x"04",x"20",x"06",x"B0",x"20",x"03",x"B5", -- 0x06C8
		x"28",x"08",x"21",x"18",x"0A",x"E5",x"CD",x"54", -- 0x06D0
		x"01",x"F1",x"3E",x"0D",x"D3",x"48",x"3E",x"00", -- 0x06D8
		x"D3",x"49",x"3E",x"0E",x"D3",x"48",x"3E",x"00", -- 0x06E0
		x"D3",x"49",x"3E",x"0F",x"D3",x"48",x"21",x"2D", -- 0x06E8
		x"02",x"39",x"7E",x"FD",x"21",x"29",x"02",x"FD", -- 0x06F0
		x"39",x"FD",x"77",x"00",x"21",x"2E",x"02",x"39", -- 0x06F8
		x"7E",x"FD",x"21",x"29",x"02",x"FD",x"39",x"FD", -- 0x0700
		x"77",x"01",x"21",x"2F",x"02",x"39",x"7E",x"FD", -- 0x0708
		x"21",x"2B",x"02",x"FD",x"39",x"FD",x"77",x"00", -- 0x0710
		x"21",x"30",x"02",x"39",x"7E",x"FD",x"21",x"2B", -- 0x0718
		x"02",x"FD",x"39",x"FD",x"77",x"01",x"FD",x"21", -- 0x0720
		x"14",x"00",x"FD",x"39",x"FD",x"36",x"00",x"00", -- 0x0728
		x"21",x"29",x"02",x"39",x"7E",x"23",x"66",x"6F", -- 0x0730
		x"FD",x"21",x"2B",x"02",x"FD",x"39",x"FD",x"5E", -- 0x0738
		x"00",x"FD",x"56",x"01",x"E5",x"D5",x"CD",x"99", -- 0x0740
		x"12",x"F1",x"F1",x"7C",x"B5",x"20",x"08",x"21", -- 0x0748
		x"37",x"0A",x"E5",x"CD",x"54",x"01",x"F1",x"21", -- 0x0750
		x"25",x"02",x"39",x"AF",x"77",x"23",x"77",x"21", -- 0x0758
		x"25",x"02",x"39",x"D5",x"FD",x"21",x"33",x"02", -- 0x0760
		x"FD",x"39",x"FD",x"E5",x"D1",x"FD",x"21",x"2F", -- 0x0768
		x"02",x"FD",x"39",x"FD",x"7E",x"00",x"86",x"12", -- 0x0770
		x"FD",x"7E",x"01",x"23",x"8E",x"13",x"12",x"D1", -- 0x0778
		x"21",x"31",x"02",x"39",x"7E",x"23",x"66",x"6F", -- 0x0780
		x"7E",x"D3",x"49",x"FD",x"21",x"25",x"02",x"FD", -- 0x0788
		x"39",x"FD",x"34",x"00",x"20",x"03",x"FD",x"34", -- 0x0790
		x"01",x"FD",x"7E",x"01",x"D6",x"02",x"38",x"BF", -- 0x0798
		x"3E",x"2E",x"F5",x"33",x"CD",x"3B",x"19",x"33", -- 0x07A0
		x"FD",x"21",x"14",x"00",x"FD",x"39",x"FD",x"34", -- 0x07A8
		x"00",x"FD",x"7E",x"00",x"D6",x"02",x"DA",x"30", -- 0x07B0
		x"07",x"21",x"19",x"09",x"E5",x"CD",x"AE",x"19", -- 0x07B8
		x"21",x"01",x"0F",x"E3",x"3E",x"0C",x"F5",x"33", -- 0x07C0
		x"CD",x"4B",x"18",x"33",x"21",x"52",x"0A",x"E3", -- 0x07C8
		x"CD",x"AE",x"19",x"F1",x"FD",x"21",x"28",x"02", -- 0x07D0
		x"FD",x"39",x"FD",x"7E",x"00",x"B7",x"20",x"08", -- 0x07D8
		x"3E",x"12",x"D3",x"48",x"3E",x"00",x"D3",x"49", -- 0x07E0
		x"21",x"FF",x"3F",x"36",x"0F",x"21",x"00",x"FF", -- 0x07E8
		x"36",x"3E",x"2E",x"01",x"36",x"F0",x"2E",x"02", -- 0x07F0
		x"36",x"D3",x"2E",x"03",x"36",x"A8",x"2E",x"04", -- 0x07F8
		x"36",x"C3",x"2E",x"05",x"36",x"00",x"2E",x"06", -- 0x0800
		x"36",x"00",x"C3",x"00",x"FF",x"21",x"35",x"02", -- 0x0808
		x"39",x"F9",x"C9",x"48",x"57",x"20",x"49",x"44", -- 0x0810
		x"20",x"3D",x"20",x"00",x"20",x"2D",x"20",x"00", -- 0x0818
		x"0A",x"0A",x"56",x"65",x"72",x"73",x"69",x"6F", -- 0x0820
		x"6E",x"20",x"00",x"0A",x"0A",x"00",x"49",x"6E", -- 0x0828
		x"69",x"74",x"69",x"61",x"6C",x"69",x"7A",x"69", -- 0x0830
		x"6E",x"67",x"20",x"53",x"44",x"20",x"43",x"61", -- 0x0838
		x"72",x"64",x"3A",x"20",x"00",x"45",x"72",x"72", -- 0x0840
		x"6F",x"72",x"20",x"6F",x"6E",x"20",x"53",x"44", -- 0x0848
		x"20",x"63",x"61",x"72",x"64",x"20",x"69",x"6E", -- 0x0850
		x"69",x"74",x"69",x"61",x"6C",x"69",x"7A",x"61", -- 0x0858
		x"74",x"69",x"6F",x"6E",x"21",x"00",x"46",x"41", -- 0x0860
		x"54",x"20",x"46",x"53",x"20",x"6E",x"6F",x"74", -- 0x0868
		x"20",x"66",x"6F",x"75",x"6E",x"64",x"21",x"00", -- 0x0870
		x"4F",x"4B",x"0A",x"0A",x"4C",x"6F",x"61",x"64", -- 0x0878
		x"69",x"6E",x"67",x"20",x"63",x"6F",x"6E",x"66", -- 0x0880
		x"69",x"67",x"20",x"66",x"69",x"6C",x"65",x"3A", -- 0x0888
		x"20",x"00",x"27",x"4D",x"53",x"58",x"31",x"46", -- 0x0890
		x"50",x"47",x"41",x"27",x"20",x"64",x"69",x"72", -- 0x0898
		x"65",x"63",x"74",x"6F",x"72",x"79",x"20",x"6E", -- 0x08A0
		x"6F",x"74",x"20",x"66",x"6F",x"75",x"6E",x"64", -- 0x08A8
		x"21",x"00",x"43",x"6F",x"6E",x"66",x"69",x"67", -- 0x08B0
		x"20",x"66",x"69",x"6C",x"65",x"20",x"6E",x"6F", -- 0x08B8
		x"74",x"20",x"66",x"6F",x"75",x"6E",x"64",x"21", -- 0x08C0
		x"00",x"43",x"6F",x"6E",x"66",x"69",x"67",x"20", -- 0x08C8
		x"66",x"69",x"6C",x"65",x"20",x"65",x"72",x"72", -- 0x08D0
		x"6F",x"72",x"21",x"00",x"45",x"72",x"72",x"6F", -- 0x08D8
		x"72",x"20",x"72",x"65",x"61",x"64",x"69",x"6E", -- 0x08E0
		x"67",x"20",x"43",x"6F",x"6E",x"66",x"69",x"67", -- 0x08E8
		x"20",x"66",x"69",x"6C",x"65",x"21",x"00",x"49", -- 0x08F0
		x"6E",x"76",x"61",x"6C",x"69",x"64",x"20",x"6B", -- 0x08F8
		x"65",x"79",x"6D",x"61",x"70",x"21",x"00",x"4F", -- 0x0900
		x"4B",x"0A",x"0A",x"5A",x"65",x"72",x"6F",x"69", -- 0x0908
		x"6E",x"67",x"20",x"52",x"41",x"4D",x"3A",x"20", -- 0x0910
		x"00",x"20",x"4F",x"4B",x"0A",x"00",x"0A",x"4C", -- 0x0918
		x"6F",x"61",x"64",x"69",x"6E",x"67",x"20",x"4D", -- 0x0920
		x"53",x"58",x"31",x"42",x"49",x"4F",x"53",x"2E", -- 0x0928
		x"52",x"4F",x"4D",x"20",x"00",x"4D",x"53",x"58", -- 0x0930
		x"31",x"42",x"49",x"4F",x"53",x"20",x"66",x"69", -- 0x0938
		x"6C",x"65",x"20",x"6E",x"6F",x"74",x"20",x"66", -- 0x0940
		x"6F",x"75",x"6E",x"64",x"21",x"00",x"4D",x"53", -- 0x0948
		x"58",x"42",x"49",x"4F",x"53",x"20",x"66",x"69", -- 0x0950
		x"6C",x"65",x"20",x"73",x"69",x"7A",x"65",x"20", -- 0x0958
		x"6D",x"75",x"73",x"74",x"20",x"62",x"65",x"20", -- 0x0960
		x"33",x"32",x"37",x"36",x"38",x"21",x"00",x"45", -- 0x0968
		x"72",x"72",x"6F",x"72",x"20",x"72",x"65",x"61", -- 0x0970
		x"64",x"69",x"6E",x"67",x"20",x"42",x"49",x"4F", -- 0x0978
		x"53",x"20",x"66",x"69",x"6C",x"65",x"21",x"00", -- 0x0980
		x"0A",x"4C",x"6F",x"61",x"64",x"69",x"6E",x"67", -- 0x0988
		x"20",x"4E",x"45",x"58",x"54",x"4F",x"52",x"2E", -- 0x0990
		x"52",x"4F",x"4D",x"20",x"00",x"4E",x"45",x"58", -- 0x0998
		x"54",x"4F",x"52",x"20",x"66",x"69",x"6C",x"65", -- 0x09A0
		x"20",x"6E",x"6F",x"74",x"20",x"66",x"6F",x"75", -- 0x09A8
		x"6E",x"64",x"21",x"00",x"4E",x"45",x"58",x"54", -- 0x09B0
		x"4F",x"52",x"20",x"66",x"69",x"6C",x"65",x"20", -- 0x09B8
		x"73",x"69",x"7A",x"65",x"20",x"6D",x"75",x"73", -- 0x09C0
		x"74",x"20",x"62",x"65",x"20",x"31",x"33",x"31", -- 0x09C8
		x"30",x"37",x"32",x"21",x"00",x"45",x"72",x"72", -- 0x09D0
		x"6F",x"72",x"20",x"72",x"65",x"61",x"64",x"69", -- 0x09D8
		x"6E",x"67",x"20",x"4E",x"45",x"58",x"54",x"4F", -- 0x09E0
		x"52",x"20",x"66",x"69",x"6C",x"65",x"21",x"00", -- 0x09E8
		x"0A",x"4C",x"6F",x"61",x"64",x"69",x"6E",x"67", -- 0x09F0
		x"20",x"4B",x"65",x"79",x"6D",x"61",x"70",x"20", -- 0x09F8
		x"00",x"4B",x"65",x"79",x"6D",x"61",x"70",x"20", -- 0x0A00
		x"66",x"69",x"6C",x"65",x"20",x"6E",x"6F",x"74", -- 0x0A08
		x"20",x"66",x"6F",x"75",x"6E",x"64",x"21",x"00", -- 0x0A10
		x"4B",x"65",x"79",x"6D",x"61",x"70",x"20",x"66", -- 0x0A18
		x"69",x"6C",x"65",x"20",x"73",x"69",x"7A",x"65", -- 0x0A20
		x"20",x"6D",x"75",x"73",x"74",x"20",x"62",x"65", -- 0x0A28
		x"20",x"31",x"30",x"32",x"34",x"21",x"00",x"45", -- 0x0A30
		x"72",x"72",x"6F",x"72",x"20",x"72",x"65",x"61", -- 0x0A38
		x"64",x"69",x"6E",x"67",x"20",x"4B",x"65",x"79", -- 0x0A40
		x"6D",x"61",x"70",x"20",x"66",x"69",x"6C",x"65", -- 0x0A48
		x"21",x"00",x"0A",x"42",x"6F",x"6F",x"74",x"69", -- 0x0A50
		x"6E",x"67",x"2E",x"2E",x"2E",x"00",x"4D",x"53", -- 0x0A58
		x"58",x"31",x"46",x"50",x"47",x"41",x"20",x"20", -- 0x0A60
		x"20",x"00",x"43",x"4F",x"4E",x"46",x"49",x"47", -- 0x0A68
		x"20",x"20",x"54",x"58",x"54",x"00",x"4E",x"45", -- 0x0A70
		x"58",x"54",x"4F",x"52",x"20",x"20",x"52",x"4F", -- 0x0A78
		x"4D",x"00",x"4D",x"53",x"58",x"31",x"42",x"49", -- 0x0A80
		x"4F",x"53",x"52",x"4F",x"4D",x"00",x"45",x"4E", -- 0x0A88
		x"20",x"20",x"20",x"20",x"20",x"20",x"4B",x"4D", -- 0x0A90
		x"50",x"00",x"50",x"54",x"42",x"52",x"20",x"20", -- 0x0A98
		x"20",x"20",x"4B",x"4D",x"50",x"00",x"46",x"52", -- 0x0AA0
		x"20",x"20",x"20",x"20",x"20",x"20",x"4B",x"4D", -- 0x0AA8
		x"50",x"00",x"53",x"50",x"41",x"20",x"20",x"20", -- 0x0AB0
		x"20",x"20",x"4B",x"4D",x"50",x"00",x"3E",x"FF", -- 0x0AB8
		x"D3",x"9E",x"06",x"0A",x"3E",x"FF",x"D3",x"9F", -- 0x0AC0
		x"10",x"FA",x"3E",x"FE",x"D3",x"9E",x"06",x"10", -- 0x0AC8
		x"3E",x"40",x"11",x"00",x"00",x"C5",x"CD",x"A6", -- 0x0AD0
		x"0B",x"C1",x"D2",x"E6",x"0A",x"10",x"F1",x"2E", -- 0x0AD8
		x"00",x"3E",x"FF",x"D3",x"9E",x"C9",x"3E",x"48", -- 0x0AE0
		x"11",x"AA",x"01",x"CD",x"B3",x"0B",x"21",x"8A", -- 0x0AE8
		x"0B",x"38",x"03",x"21",x"98",x"0B",x"01",x"78", -- 0x0AF0
		x"00",x"C5",x"CD",x"0D",x"0B",x"C1",x"D2",x"0E", -- 0x0AF8
		x"0B",x"10",x"F6",x"0D",x"20",x"F3",x"2E",x"00", -- 0x0B00
		x"3E",x"FF",x"D3",x"9E",x"C9",x"E9",x"3E",x"7A", -- 0x0B08
		x"11",x"00",x"00",x"CD",x"B3",x"0B",x"DA",x"06", -- 0x0B10
		x"0B",x"78",x"E6",x"40",x"32",x"00",x"40",x"CC", -- 0x0B18
		x"31",x"0B",x"3E",x"FF",x"D3",x"9E",x"3A",x"00", -- 0x0B20
		x"40",x"2E",x"03",x"FE",x"40",x"C8",x"2E",x"02", -- 0x0B28
		x"C9",x"3E",x"50",x"01",x"00",x"00",x"11",x"00", -- 0x0B30
		x"02",x"C3",x"91",x"0B",x"FD",x"21",x"00",x"00", -- 0x0B38
		x"FD",x"39",x"FD",x"5E",x"02",x"FD",x"56",x"03", -- 0x0B40
		x"FD",x"4E",x"04",x"FD",x"46",x"05",x"FD",x"6E", -- 0x0B48
		x"06",x"FD",x"66",x"07",x"3E",x"FE",x"D3",x"9E", -- 0x0B50
		x"3A",x"00",x"40",x"B7",x"CC",x"7E",x"0B",x"3E", -- 0x0B58
		x"51",x"CD",x"91",x"0B",x"30",x"03",x"2E",x"00", -- 0x0B60
		x"C9",x"CD",x"F3",x"0B",x"38",x"F8",x"01",x"9F", -- 0x0B68
		x"00",x"ED",x"B2",x"ED",x"B2",x"00",x"DB",x"9F", -- 0x0B70
		x"00",x"DB",x"9F",x"2E",x"01",x"C9",x"41",x"4A", -- 0x0B78
		x"53",x"1E",x"00",x"CB",x"22",x"CB",x"11",x"CB", -- 0x0B80
		x"10",x"C9",x"3E",x"41",x"01",x"00",x"00",x"50", -- 0x0B88
		x"59",x"CD",x"CC",x"0B",x"B7",x"C8",x"37",x"C9", -- 0x0B90
		x"3E",x"77",x"CD",x"8C",x"0B",x"3E",x"69",x"01", -- 0x0B98
		x"00",x"40",x"51",x"59",x"18",x"EB",x"01",x"00", -- 0x0BA0
		x"00",x"CD",x"CC",x"0B",x"47",x"E6",x"FE",x"78", -- 0x0BA8
		x"20",x"E4",x"C9",x"CD",x"A6",x"0B",x"D8",x"F5", -- 0x0BB0
		x"CD",x"01",x"0C",x"67",x"CD",x"01",x"0C",x"6F", -- 0x0BB8
		x"CD",x"01",x"0C",x"57",x"CD",x"01",x"0C",x"5F", -- 0x0BC0
		x"44",x"4D",x"F1",x"C9",x"D3",x"9F",x"F5",x"78", -- 0x0BC8
		x"00",x"D3",x"9F",x"79",x"00",x"D3",x"9F",x"7A", -- 0x0BD0
		x"00",x"D3",x"9F",x"7B",x"00",x"D3",x"9F",x"F1", -- 0x0BD8
		x"FE",x"40",x"06",x"95",x"28",x"08",x"FE",x"48", -- 0x0BE0
		x"06",x"87",x"28",x"02",x"06",x"FF",x"78",x"D3", -- 0x0BE8
		x"9F",x"18",x"0E",x"06",x"0A",x"C5",x"CD",x"01", -- 0x0BF0
		x"0C",x"C1",x"FE",x"FE",x"C8",x"10",x"F6",x"37", -- 0x0BF8
		x"C9",x"01",x"64",x"00",x"DB",x"9F",x"FE",x"FF", -- 0x0C00
		x"C0",x"10",x"F9",x"0D",x"20",x"F6",x"C9",x"C1", -- 0x0C08
		x"E1",x"E5",x"C5",x"46",x"23",x"4E",x"23",x"5E", -- 0x0C10
		x"23",x"56",x"68",x"61",x"C9",x"C1",x"E1",x"E5", -- 0x0C18
		x"C5",x"7E",x"23",x"66",x"6F",x"C9",x"F5",x"F5", -- 0x0C20
		x"21",x"06",x"00",x"39",x"5E",x"23",x"56",x"21", -- 0x0C28
		x"08",x"00",x"39",x"7E",x"FD",x"21",x"00",x"00", -- 0x0C30
		x"FD",x"39",x"FD",x"77",x"00",x"21",x"09",x"00", -- 0x0C38
		x"39",x"7E",x"FD",x"21",x"00",x"00",x"FD",x"39", -- 0x0C40
		x"FD",x"77",x"01",x"01",x"00",x"00",x"21",x"0A", -- 0x0C48
		x"00",x"39",x"79",x"96",x"78",x"23",x"9E",x"E2", -- 0x0C50
		x"5C",x"0C",x"EE",x"80",x"F2",x"9C",x"0C",x"1A", -- 0x0C58
		x"FD",x"21",x"03",x"00",x"FD",x"39",x"FD",x"77", -- 0x0C60
		x"00",x"13",x"E1",x"E5",x"7E",x"FD",x"21",x"02", -- 0x0C68
		x"00",x"FD",x"39",x"FD",x"77",x"00",x"FD",x"21", -- 0x0C70
		x"00",x"00",x"FD",x"39",x"FD",x"34",x"00",x"20", -- 0x0C78
		x"03",x"FD",x"34",x"01",x"21",x"03",x"00",x"39", -- 0x0C80
		x"7E",x"FD",x"21",x"02",x"00",x"FD",x"39",x"FD", -- 0x0C88
		x"96",x"00",x"28",x"05",x"21",x"00",x"00",x"18", -- 0x0C90
		x"06",x"03",x"18",x"B2",x"21",x"01",x"00",x"F1", -- 0x0C98
		x"F1",x"C9",x"ED",x"5B",x"02",x"40",x"ED",x"4B", -- 0x0CA0
		x"04",x"40",x"21",x"02",x"00",x"39",x"7E",x"83", -- 0x0CA8
		x"77",x"23",x"7E",x"8A",x"77",x"23",x"7E",x"89", -- 0x0CB0
		x"77",x"23",x"7E",x"88",x"77",x"ED",x"5B",x"0E", -- 0x0CB8
		x"40",x"ED",x"4B",x"10",x"40",x"FD",x"21",x"02", -- 0x0CC0
		x"00",x"FD",x"39",x"FD",x"7E",x"00",x"93",x"20", -- 0x0CC8
		x"16",x"FD",x"7E",x"01",x"92",x"20",x"10",x"FD", -- 0x0CD0
		x"7E",x"02",x"91",x"20",x"0A",x"FD",x"7E",x"03", -- 0x0CD8
		x"90",x"20",x"04",x"21",x"01",x"00",x"C9",x"21", -- 0x0CE0
		x"24",x"40",x"E5",x"FD",x"21",x"04",x"00",x"FD", -- 0x0CE8
		x"39",x"FD",x"6E",x"02",x"FD",x"66",x"03",x"E5", -- 0x0CF0
		x"FD",x"6E",x"00",x"FD",x"66",x"01",x"E5",x"CD", -- 0x0CF8
		x"3C",x"0B",x"F1",x"F1",x"F1",x"7D",x"B7",x"28", -- 0x0D00
		x"10",x"11",x"0E",x"40",x"21",x"02",x"00",x"39", -- 0x0D08
		x"01",x"04",x"00",x"ED",x"B0",x"21",x"01",x"00", -- 0x0D10
		x"C9",x"21",x"00",x"00",x"C9",x"F5",x"F5",x"F5", -- 0x0D18
		x"F5",x"11",x"06",x"40",x"21",x"04",x"00",x"39", -- 0x0D20
		x"EB",x"01",x"04",x"00",x"ED",x"B0",x"FD",x"21", -- 0x0D28
		x"0A",x"00",x"FD",x"39",x"FD",x"7E",x"00",x"C6", -- 0x0D30
		x"FE",x"5F",x"FD",x"7E",x"01",x"CE",x"FF",x"57", -- 0x0D38
		x"FD",x"7E",x"02",x"CE",x"FF",x"4F",x"FD",x"7E", -- 0x0D40
		x"03",x"CE",x"FF",x"47",x"3A",x"01",x"40",x"FD", -- 0x0D48
		x"21",x"00",x"00",x"FD",x"39",x"FD",x"77",x"00", -- 0x0D50
		x"FD",x"36",x"01",x"00",x"FD",x"36",x"02",x"00", -- 0x0D58
		x"FD",x"36",x"03",x"00",x"FD",x"6E",x"02",x"FD", -- 0x0D60
		x"66",x"03",x"E5",x"FD",x"6E",x"00",x"FD",x"66", -- 0x0D68
		x"01",x"E5",x"C5",x"D5",x"CD",x"EC",x"19",x"F1", -- 0x0D70
		x"F1",x"F1",x"F1",x"4D",x"44",x"FD",x"21",x"04", -- 0x0D78
		x"00",x"FD",x"39",x"FD",x"7E",x"00",x"81",x"4F", -- 0x0D80
		x"FD",x"7E",x"01",x"88",x"47",x"FD",x"7E",x"02", -- 0x0D88
		x"8B",x"5F",x"FD",x"7E",x"03",x"8A",x"57",x"69", -- 0x0D90
		x"60",x"F1",x"F1",x"F1",x"F1",x"C9",x"F5",x"FD", -- 0x0D98
		x"21",x"04",x"00",x"FD",x"39",x"FD",x"6E",x"00", -- 0x0DA0
		x"FD",x"66",x"01",x"FD",x"5E",x"02",x"FD",x"56", -- 0x0DA8
		x"03",x"F1",x"06",x"08",x"CB",x"3A",x"CB",x"1B", -- 0x0DB0
		x"CB",x"1C",x"CB",x"1D",x"10",x"F6",x"D5",x"E5", -- 0x0DB8
		x"CD",x"A2",x"0C",x"F1",x"F1",x"4D",x"7C",x"B1", -- 0x0DC0
		x"20",x"06",x"21",x"00",x"00",x"5D",x"54",x"C9", -- 0x0DC8
		x"11",x"24",x"40",x"FD",x"21",x"02",x"00",x"FD", -- 0x0DD0
		x"39",x"FD",x"6E",x"00",x"26",x"00",x"01",x"00", -- 0x0DD8
		x"00",x"29",x"CB",x"11",x"CB",x"10",x"19",x"E5", -- 0x0DE0
		x"CD",x"1D",x"0C",x"F1",x"11",x"00",x"00",x"C9", -- 0x0DE8
		x"FD",x"21",x"02",x"00",x"FD",x"39",x"FD",x"7E", -- 0x0DF0
		x"00",x"E6",x"F8",x"6F",x"FD",x"66",x"01",x"11", -- 0x0DF8
		x"00",x"00",x"7D",x"D6",x"F8",x"20",x"0E",x"24", -- 0x0E00
		x"20",x"0B",x"7B",x"B7",x"20",x"07",x"B2",x"20", -- 0x0E08
		x"04",x"3E",x"01",x"18",x"01",x"AF",x"6F",x"17", -- 0x0E10
		x"9F",x"67",x"C9",x"F5",x"F5",x"F5",x"F5",x"3A", -- 0x0E18
		x"34",x"42",x"33",x"F5",x"33",x"21",x"3A",x"42", -- 0x0E20
		x"E5",x"CD",x"1D",x"0C",x"F1",x"FD",x"21",x"01", -- 0x0E28
		x"00",x"FD",x"39",x"FD",x"75",x"00",x"FD",x"74", -- 0x0E30
		x"01",x"21",x"00",x"00",x"22",x"12",x"40",x"22", -- 0x0E38
		x"14",x"40",x"ED",x"5B",x"02",x"40",x"ED",x"4B", -- 0x0E40
		x"04",x"40",x"ED",x"53",x"16",x"40",x"ED",x"43", -- 0x0E48
		x"18",x"40",x"21",x"00",x"00",x"39",x"7E",x"FD", -- 0x0E50
		x"21",x"03",x"00",x"FD",x"39",x"FD",x"77",x"00", -- 0x0E58
		x"FD",x"21",x"03",x"00",x"FD",x"39",x"FD",x"7E", -- 0x0E60
		x"00",x"B7",x"28",x"44",x"11",x"16",x"40",x"21", -- 0x0E68
		x"04",x"00",x"39",x"EB",x"01",x"04",x"00",x"ED", -- 0x0E70
		x"B0",x"21",x"01",x"00",x"39",x"5E",x"23",x"56", -- 0x0E78
		x"01",x"00",x"00",x"FD",x"21",x"04",x"00",x"FD", -- 0x0E80
		x"39",x"FD",x"7E",x"00",x"83",x"5F",x"FD",x"7E", -- 0x0E88
		x"01",x"8A",x"57",x"FD",x"7E",x"02",x"89",x"4F", -- 0x0E90
		x"FD",x"7E",x"03",x"88",x"47",x"ED",x"53",x"16", -- 0x0E98
		x"40",x"ED",x"43",x"18",x"40",x"FD",x"21",x"03", -- 0x0EA0
		x"00",x"FD",x"39",x"FD",x"35",x"00",x"18",x"B0", -- 0x0EA8
		x"21",x"35",x"42",x"E5",x"CD",x"1D",x"0C",x"F1", -- 0x0EB0
		x"EB",x"06",x"04",x"CB",x"3A",x"CB",x"1B",x"10", -- 0x0EB8
		x"FA",x"ED",x"53",x"1A",x"40",x"D5",x"11",x"16", -- 0x0EC0
		x"40",x"21",x"06",x"00",x"39",x"EB",x"01",x"04", -- 0x0EC8
		x"00",x"ED",x"B0",x"D1",x"01",x"00",x"00",x"FD", -- 0x0ED0
		x"21",x"04",x"00",x"FD",x"39",x"FD",x"7E",x"00", -- 0x0ED8
		x"83",x"5F",x"FD",x"7E",x"01",x"8A",x"57",x"FD", -- 0x0EE0
		x"7E",x"02",x"89",x"4F",x"FD",x"7E",x"03",x"88", -- 0x0EE8
		x"47",x"ED",x"53",x"06",x"40",x"ED",x"43",x"08", -- 0x0EF0
		x"40",x"21",x"00",x"00",x"22",x"1C",x"40",x"22", -- 0x0EF8
		x"1E",x"40",x"ED",x"5B",x"16",x"40",x"ED",x"4B", -- 0x0F00
		x"18",x"40",x"ED",x"53",x"20",x"40",x"ED",x"43", -- 0x0F08
		x"22",x"40",x"F1",x"F1",x"F1",x"F1",x"C9",x"F5", -- 0x0F10
		x"F5",x"21",x"24",x"42",x"E5",x"21",x"00",x"00", -- 0x0F18
		x"E5",x"21",x"00",x"00",x"E5",x"CD",x"3C",x"0B", -- 0x0F20
		x"F1",x"F1",x"F1",x"7D",x"B7",x"20",x"06",x"21", -- 0x0F28
		x"00",x"00",x"C3",x"22",x"10",x"3A",x"22",x"44", -- 0x0F30
		x"D6",x"55",x"20",x"07",x"3A",x"23",x"44",x"D6", -- 0x0F38
		x"AA",x"28",x"06",x"21",x"00",x"00",x"C3",x"22", -- 0x0F40
		x"10",x"3A",x"E6",x"43",x"FE",x"04",x"28",x"04", -- 0x0F48
		x"D6",x"06",x"20",x"04",x"0E",x"01",x"18",x"10", -- 0x0F50
		x"3A",x"5D",x"42",x"D6",x"31",x"20",x"03",x"4F", -- 0x0F58
		x"18",x"06",x"21",x"00",x"00",x"C3",x"22",x"10", -- 0x0F60
		x"79",x"B7",x"28",x"1C",x"21",x"EA",x"43",x"E5", -- 0x0F68
		x"CD",x"0F",x"0C",x"F1",x"FD",x"21",x"00",x"00", -- 0x0F70
		x"FD",x"39",x"FD",x"75",x"00",x"FD",x"74",x"01", -- 0x0F78
		x"FD",x"73",x"02",x"FD",x"72",x"03",x"18",x"13", -- 0x0F80
		x"AF",x"FD",x"21",x"00",x"00",x"FD",x"39",x"FD", -- 0x0F88
		x"77",x"00",x"FD",x"77",x"01",x"FD",x"77",x"02", -- 0x0F90
		x"FD",x"77",x"03",x"21",x"24",x"42",x"E5",x"FD", -- 0x0F98
		x"21",x"02",x"00",x"FD",x"39",x"FD",x"6E",x"02", -- 0x0FA0
		x"FD",x"66",x"03",x"E5",x"FD",x"6E",x"00",x"FD", -- 0x0FA8
		x"66",x"01",x"E5",x"CD",x"3C",x"0B",x"F1",x"F1", -- 0x0FB0
		x"F1",x"7D",x"B7",x"20",x"05",x"21",x"00",x"00", -- 0x0FB8
		x"18",x"60",x"3A",x"22",x"44",x"D6",x"55",x"20", -- 0x0FC0
		x"07",x"3A",x"23",x"44",x"D6",x"AA",x"28",x"05", -- 0x0FC8
		x"21",x"00",x"00",x"18",x"4D",x"3A",x"2F",x"42", -- 0x0FD0
		x"B7",x"20",x"07",x"3A",x"30",x"42",x"D6",x"02", -- 0x0FD8
		x"28",x"05",x"21",x"00",x"00",x"18",x"3B",x"11", -- 0x0FE0
		x"01",x"40",x"3A",x"31",x"42",x"12",x"21",x"32", -- 0x0FE8
		x"42",x"E5",x"CD",x"1D",x"0C",x"F1",x"EB",x"01", -- 0x0FF0
		x"00",x"00",x"FD",x"21",x"00",x"00",x"FD",x"39", -- 0x0FF8
		x"FD",x"7E",x"00",x"83",x"5F",x"FD",x"7E",x"01", -- 0x1000
		x"8A",x"57",x"FD",x"7E",x"02",x"89",x"4F",x"FD", -- 0x1008
		x"7E",x"03",x"88",x"47",x"ED",x"53",x"02",x"40", -- 0x1010
		x"ED",x"43",x"04",x"40",x"CD",x"1B",x"0E",x"21", -- 0x1018
		x"01",x"00",x"F1",x"F1",x"C9",x"21",x"EA",x"FF", -- 0x1020
		x"39",x"F9",x"11",x"20",x"40",x"21",x"12",x"00", -- 0x1028
		x"39",x"EB",x"01",x"04",x"00",x"ED",x"B0",x"2A", -- 0x1030
		x"1A",x"40",x"FD",x"21",x"05",x"00",x"FD",x"39", -- 0x1038
		x"FD",x"75",x"00",x"21",x"05",x"00",x"39",x"7E", -- 0x1040
		x"B7",x"CA",x"30",x"12",x"21",x"24",x"42",x"E5", -- 0x1048
		x"FD",x"21",x"14",x"00",x"FD",x"39",x"FD",x"6E", -- 0x1050
		x"02",x"FD",x"66",x"03",x"E5",x"FD",x"6E",x"00", -- 0x1058
		x"FD",x"66",x"01",x"E5",x"CD",x"3C",x"0B",x"F1", -- 0x1060
		x"F1",x"F1",x"7D",x"B7",x"20",x"06",x"21",x"00", -- 0x1068
		x"00",x"C3",x"33",x"12",x"FD",x"21",x"00",x"00", -- 0x1070
		x"FD",x"39",x"FD",x"36",x"00",x"24",x"FD",x"36", -- 0x1078
		x"01",x"42",x"FD",x"7E",x"00",x"FD",x"21",x"03", -- 0x1080
		x"00",x"FD",x"39",x"FD",x"77",x"00",x"21",x"01", -- 0x1088
		x"00",x"39",x"7E",x"FD",x"21",x"03",x"00",x"FD", -- 0x1090
		x"39",x"FD",x"77",x"01",x"FD",x"21",x"02",x"00", -- 0x1098
		x"FD",x"39",x"FD",x"36",x"00",x"00",x"FD",x"21", -- 0x10A0
		x"03",x"00",x"FD",x"39",x"FD",x"6E",x"00",x"FD", -- 0x10A8
		x"66",x"01",x"7E",x"FE",x"E5",x"CA",x"D2",x"11", -- 0x10B0
		x"B7",x"CA",x"D2",x"11",x"FD",x"6E",x"00",x"FD", -- 0x10B8
		x"66",x"01",x"01",x"0B",x"00",x"C5",x"FD",x"21", -- 0x10C0
		x"1C",x"00",x"FD",x"39",x"FD",x"4E",x"00",x"FD", -- 0x10C8
		x"46",x"01",x"C5",x"E5",x"CD",x"26",x"0C",x"F1", -- 0x10D0
		x"F1",x"F1",x"7C",x"B5",x"CA",x"D2",x"11",x"21", -- 0x10D8
		x"18",x"00",x"39",x"7E",x"FD",x"21",x"0E",x"00", -- 0x10E0
		x"FD",x"39",x"FD",x"77",x"00",x"21",x"19",x"00", -- 0x10E8
		x"39",x"7E",x"FD",x"21",x"0E",x"00",x"FD",x"39", -- 0x10F0
		x"FD",x"77",x"01",x"E1",x"E5",x"11",x"0B",x"00", -- 0x10F8
		x"19",x"7E",x"FD",x"6E",x"00",x"FD",x"66",x"01", -- 0x1100
		x"77",x"21",x"10",x"00",x"39",x"FD",x"7E",x"00", -- 0x1108
		x"C6",x"01",x"77",x"FD",x"7E",x"01",x"CE",x"00", -- 0x1110
		x"23",x"77",x"FD",x"21",x"00",x"00",x"FD",x"39", -- 0x1118
		x"FD",x"7E",x"00",x"C6",x"1C",x"5F",x"FD",x"7E", -- 0x1120
		x"01",x"CE",x"00",x"57",x"D5",x"CD",x"0F",x"0C", -- 0x1128
		x"F1",x"FD",x"21",x"0A",x"00",x"FD",x"39",x"FD", -- 0x1130
		x"72",x"03",x"FD",x"73",x"02",x"FD",x"74",x"01", -- 0x1138
		x"FD",x"75",x"00",x"21",x"10",x"00",x"39",x"5E", -- 0x1140
		x"23",x"56",x"21",x"0A",x"00",x"39",x"01",x"04", -- 0x1148
		x"00",x"ED",x"B0",x"21",x"0A",x"00",x"39",x"FD", -- 0x1150
		x"21",x"0E",x"00",x"FD",x"39",x"FD",x"7E",x"00", -- 0x1158
		x"C6",x"05",x"77",x"FD",x"7E",x"01",x"CE",x"00", -- 0x1160
		x"23",x"77",x"21",x"10",x"00",x"39",x"FD",x"21", -- 0x1168
		x"00",x"00",x"FD",x"39",x"FD",x"7E",x"00",x"C6", -- 0x1170
		x"1A",x"77",x"FD",x"7E",x"01",x"CE",x"00",x"23", -- 0x1178
		x"77",x"21",x"10",x"00",x"39",x"4E",x"23",x"46", -- 0x1180
		x"C5",x"CD",x"1D",x"0C",x"F1",x"FD",x"21",x"10", -- 0x1188
		x"00",x"FD",x"39",x"FD",x"74",x"01",x"FD",x"75", -- 0x1190
		x"00",x"21",x"10",x"00",x"39",x"7E",x"FD",x"21", -- 0x1198
		x"06",x"00",x"FD",x"39",x"FD",x"77",x"00",x"21", -- 0x11A0
		x"11",x"00",x"39",x"7E",x"FD",x"21",x"06",x"00", -- 0x11A8
		x"FD",x"39",x"FD",x"77",x"01",x"FD",x"36",x"02", -- 0x11B0
		x"00",x"FD",x"36",x"03",x"00",x"21",x"0A",x"00", -- 0x11B8
		x"39",x"5E",x"23",x"56",x"21",x"06",x"00",x"39", -- 0x11C0
		x"01",x"04",x"00",x"ED",x"B0",x"21",x"01",x"00", -- 0x11C8
		x"18",x"61",x"21",x"03",x"00",x"39",x"7E",x"C6", -- 0x11D0
		x"20",x"77",x"23",x"7E",x"CE",x"00",x"77",x"21", -- 0x11D8
		x"03",x"00",x"39",x"7E",x"FD",x"21",x"00",x"00", -- 0x11E0
		x"FD",x"39",x"FD",x"77",x"00",x"21",x"04",x"00", -- 0x11E8
		x"39",x"7E",x"FD",x"21",x"00",x"00",x"FD",x"39", -- 0x11F0
		x"FD",x"77",x"01",x"FD",x"21",x"02",x"00",x"FD", -- 0x11F8
		x"39",x"FD",x"34",x"00",x"FD",x"7E",x"00",x"D6", -- 0x1200
		x"10",x"DA",x"A6",x"10",x"FD",x"21",x"12",x"00", -- 0x1208
		x"FD",x"39",x"FD",x"34",x"00",x"20",x"0D",x"FD", -- 0x1210
		x"34",x"01",x"20",x"08",x"FD",x"34",x"02",x"20", -- 0x1218
		x"03",x"FD",x"34",x"03",x"FD",x"21",x"05",x"00", -- 0x1220
		x"FD",x"39",x"FD",x"35",x"00",x"C3",x"43",x"10", -- 0x1228
		x"21",x"00",x"00",x"FD",x"21",x"16",x"00",x"FD", -- 0x1230
		x"39",x"FD",x"F9",x"C9",x"F5",x"21",x"06",x"00", -- 0x1238
		x"39",x"4E",x"23",x"46",x"C5",x"21",x"06",x"00", -- 0x1240
		x"39",x"4E",x"23",x"46",x"C5",x"CD",x"25",x"10", -- 0x1248
		x"F1",x"F1",x"7C",x"B5",x"20",x"05",x"21",x"00", -- 0x1250
		x"00",x"18",x"3C",x"FD",x"21",x"04",x"00",x"FD", -- 0x1258
		x"39",x"FD",x"5E",x"00",x"FD",x"56",x"01",x"1A", -- 0x1260
		x"E6",x"18",x"28",x"05",x"21",x"00",x"00",x"18", -- 0x1268
		x"26",x"21",x"09",x"00",x"19",x"E3",x"EB",x"11", -- 0x1270
		x"05",x"00",x"19",x"5E",x"23",x"56",x"23",x"4E", -- 0x1278
		x"23",x"46",x"C5",x"D5",x"CD",x"1D",x"0D",x"F1", -- 0x1280
		x"F1",x"4D",x"44",x"E1",x"E5",x"71",x"23",x"70", -- 0x1288
		x"23",x"73",x"23",x"72",x"21",x"01",x"00",x"F1", -- 0x1290
		x"C9",x"F5",x"F5",x"F5",x"F5",x"21",x"0A",x"00", -- 0x1298
		x"39",x"5E",x"23",x"56",x"21",x"09",x"00",x"19", -- 0x12A0
		x"FD",x"21",x"06",x"00",x"FD",x"39",x"FD",x"75", -- 0x12A8
		x"00",x"FD",x"74",x"01",x"D5",x"FD",x"5E",x"00", -- 0x12B0
		x"FD",x"56",x"01",x"21",x"04",x"00",x"39",x"EB", -- 0x12B8
		x"01",x"04",x"00",x"ED",x"B0",x"D1",x"21",x"05", -- 0x12C0
		x"00",x"19",x"E3",x"E1",x"E5",x"5E",x"23",x"56", -- 0x12C8
		x"23",x"4E",x"23",x"46",x"1C",x"20",x"07",x"14", -- 0x12D0
		x"20",x"04",x"0C",x"20",x"01",x"04",x"C5",x"D5", -- 0x12D8
		x"CD",x"1D",x"0D",x"F1",x"F1",x"4D",x"44",x"FD", -- 0x12E0
		x"21",x"02",x"00",x"FD",x"39",x"FD",x"7E",x"00", -- 0x12E8
		x"91",x"20",x"5E",x"FD",x"7E",x"01",x"90",x"20", -- 0x12F0
		x"58",x"FD",x"7E",x"02",x"93",x"20",x"52",x"FD", -- 0x12F8
		x"7E",x"03",x"92",x"20",x"4C",x"E1",x"E5",x"5E", -- 0x1300
		x"23",x"56",x"23",x"4E",x"23",x"46",x"C5",x"D5", -- 0x1308
		x"CD",x"9E",x"0D",x"F1",x"F1",x"4D",x"44",x"E1", -- 0x1310
		x"E5",x"71",x"23",x"70",x"23",x"73",x"23",x"72", -- 0x1318
		x"D5",x"C5",x"CD",x"F0",x"0D",x"F1",x"F1",x"7C", -- 0x1320
		x"B5",x"28",x"05",x"21",x"FF",x"FF",x"18",x"71", -- 0x1328
		x"E1",x"E5",x"5E",x"23",x"56",x"23",x"4E",x"23", -- 0x1330
		x"46",x"C5",x"D5",x"CD",x"1D",x"0D",x"F1",x"F1", -- 0x1338
		x"4D",x"44",x"21",x"06",x"00",x"39",x"7E",x"23", -- 0x1340
		x"66",x"6F",x"71",x"23",x"70",x"23",x"73",x"23", -- 0x1348
		x"72",x"FD",x"21",x"06",x"00",x"FD",x"39",x"FD", -- 0x1350
		x"6E",x"00",x"FD",x"66",x"01",x"5E",x"23",x"56", -- 0x1358
		x"23",x"4E",x"23",x"46",x"7B",x"21",x"02",x"00", -- 0x1360
		x"39",x"C6",x"01",x"77",x"7A",x"CE",x"00",x"23", -- 0x1368
		x"77",x"79",x"CE",x"00",x"23",x"77",x"78",x"CE", -- 0x1370
		x"00",x"23",x"77",x"D5",x"C5",x"FD",x"5E",x"00", -- 0x1378
		x"FD",x"56",x"01",x"21",x"06",x"00",x"39",x"01", -- 0x1380
		x"04",x"00",x"ED",x"B0",x"C1",x"D1",x"21",x"0C", -- 0x1388
		x"00",x"39",x"7E",x"23",x"66",x"6F",x"E5",x"C5", -- 0x1390
		x"D5",x"CD",x"3C",x"0B",x"F1",x"F1",x"F1",x"26", -- 0x1398
		x"00",x"F1",x"F1",x"F1",x"F1",x"C9",x"21",x"EF", -- 0x13A0
		x"FF",x"39",x"F9",x"21",x"00",x"00",x"39",x"5D", -- 0x13A8
		x"54",x"D5",x"FD",x"21",x"15",x"00",x"FD",x"39", -- 0x13B0
		x"FD",x"4E",x"00",x"FD",x"46",x"01",x"C5",x"E5", -- 0x13B8
		x"CD",x"25",x"10",x"F1",x"F1",x"D1",x"7C",x"B5", -- 0x13C0
		x"20",x"05",x"21",x"00",x"00",x"18",x"42",x"1A", -- 0x13C8
		x"CB",x"67",x"20",x"05",x"21",x"00",x"00",x"18", -- 0x13D0
		x"38",x"13",x"13",x"13",x"13",x"13",x"D5",x"21", -- 0x13D8
		x"0F",x"00",x"39",x"EB",x"01",x"04",x"00",x"ED", -- 0x13E0
		x"B0",x"11",x"1C",x"40",x"21",x"0F",x"00",x"39", -- 0x13E8
		x"01",x"04",x"00",x"ED",x"B0",x"E1",x"5E",x"23", -- 0x13F0
		x"56",x"23",x"4E",x"23",x"46",x"C5",x"D5",x"CD", -- 0x13F8
		x"1D",x"0D",x"F1",x"F1",x"4D",x"44",x"ED",x"43", -- 0x1400
		x"20",x"40",x"ED",x"53",x"22",x"40",x"21",x"01", -- 0x1408
		x"00",x"FD",x"21",x"11",x"00",x"FD",x"39",x"FD", -- 0x1410
		x"F9",x"C9",x"21",x"03",x"00",x"39",x"7E",x"D3", -- 0x1418
		x"99",x"21",x"02",x"00",x"39",x"7E",x"E6",x"07", -- 0x1420
		x"CB",x"FF",x"D3",x"99",x"C9",x"28",x"00",x"00", -- 0x1428
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10", -- 0x1430
		x"10",x"10",x"10",x"00",x"10",x"00",x"00",x"24", -- 0x1438
		x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24", -- 0x1440
		x"7E",x"24",x"24",x"7E",x"24",x"00",x"00",x"08", -- 0x1448
		x"3E",x"28",x"3E",x"0A",x"3E",x"08",x"00",x"62", -- 0x1450
		x"64",x"08",x"10",x"26",x"46",x"00",x"00",x"10", -- 0x1458
		x"28",x"10",x"2A",x"44",x"3A",x"00",x"00",x"08", -- 0x1460
		x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"04", -- 0x1468
		x"08",x"08",x"08",x"08",x"04",x"00",x"00",x"20", -- 0x1470
		x"10",x"10",x"10",x"10",x"20",x"00",x"00",x"00", -- 0x1478
		x"14",x"08",x"3E",x"08",x"14",x"00",x"00",x"00", -- 0x1480
		x"08",x"08",x"3E",x"08",x"08",x"00",x"00",x"00", -- 0x1488
		x"00",x"00",x"00",x"08",x"08",x"10",x"00",x"00", -- 0x1490
		x"00",x"00",x"3E",x"00",x"00",x"00",x"00",x"00", -- 0x1498
		x"00",x"00",x"00",x"18",x"18",x"00",x"00",x"00", -- 0x14A0
		x"02",x"04",x"08",x"10",x"20",x"00",x"00",x"3C", -- 0x14A8
		x"46",x"4A",x"52",x"62",x"3C",x"00",x"00",x"18", -- 0x14B0
		x"28",x"08",x"08",x"08",x"3E",x"00",x"00",x"3C", -- 0x14B8
		x"42",x"02",x"3C",x"40",x"7E",x"00",x"00",x"3C", -- 0x14C0
		x"42",x"0C",x"02",x"42",x"3C",x"00",x"00",x"08", -- 0x14C8
		x"18",x"28",x"48",x"7E",x"08",x"00",x"00",x"7E", -- 0x14D0
		x"40",x"7C",x"02",x"42",x"3C",x"00",x"00",x"3C", -- 0x14D8
		x"40",x"7C",x"42",x"42",x"3C",x"00",x"00",x"7E", -- 0x14E0
		x"02",x"04",x"08",x"10",x"10",x"00",x"00",x"3C", -- 0x14E8
		x"42",x"3C",x"42",x"42",x"3C",x"00",x"00",x"3C", -- 0x14F0
		x"42",x"42",x"3E",x"02",x"3C",x"00",x"00",x"00", -- 0x14F8
		x"00",x"10",x"00",x"00",x"10",x"00",x"00",x"00", -- 0x1500
		x"10",x"00",x"00",x"10",x"10",x"20",x"00",x"00", -- 0x1508
		x"04",x"08",x"10",x"08",x"04",x"00",x"00",x"00", -- 0x1510
		x"00",x"3E",x"00",x"3E",x"00",x"00",x"00",x"00", -- 0x1518
		x"20",x"10",x"08",x"10",x"20",x"00",x"00",x"3C", -- 0x1520
		x"42",x"04",x"08",x"00",x"08",x"00",x"00",x"3C", -- 0x1528
		x"4A",x"56",x"5E",x"40",x"3C",x"00",x"00",x"3C", -- 0x1530
		x"42",x"42",x"7E",x"42",x"42",x"00",x"00",x"7C", -- 0x1538
		x"42",x"7C",x"42",x"42",x"7C",x"00",x"00",x"3C", -- 0x1540
		x"42",x"40",x"40",x"42",x"3C",x"00",x"00",x"78", -- 0x1548
		x"44",x"42",x"42",x"44",x"78",x"00",x"00",x"7E", -- 0x1550
		x"40",x"7C",x"40",x"40",x"7E",x"00",x"00",x"7E", -- 0x1558
		x"40",x"7C",x"40",x"40",x"40",x"00",x"00",x"3C", -- 0x1560
		x"42",x"40",x"4E",x"42",x"3C",x"00",x"00",x"42", -- 0x1568
		x"42",x"7E",x"42",x"42",x"42",x"00",x"00",x"3E", -- 0x1570
		x"08",x"08",x"08",x"08",x"3E",x"00",x"00",x"02", -- 0x1578
		x"02",x"02",x"42",x"42",x"3C",x"00",x"00",x"44", -- 0x1580
		x"48",x"70",x"48",x"44",x"42",x"00",x"00",x"40", -- 0x1588
		x"40",x"40",x"40",x"40",x"7E",x"00",x"00",x"42", -- 0x1590
		x"66",x"5A",x"42",x"42",x"42",x"00",x"00",x"42", -- 0x1598
		x"62",x"52",x"4A",x"46",x"42",x"00",x"00",x"3C", -- 0x15A0
		x"42",x"42",x"42",x"42",x"3C",x"00",x"00",x"7C", -- 0x15A8
		x"42",x"42",x"7C",x"40",x"40",x"00",x"00",x"3C", -- 0x15B0
		x"42",x"42",x"52",x"4A",x"3C",x"00",x"00",x"7C", -- 0x15B8
		x"42",x"42",x"7C",x"44",x"42",x"00",x"00",x"3C", -- 0x15C0
		x"40",x"3C",x"02",x"42",x"3C",x"00",x"00",x"FE", -- 0x15C8
		x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"42", -- 0x15D0
		x"42",x"42",x"42",x"42",x"3C",x"00",x"00",x"42", -- 0x15D8
		x"42",x"42",x"42",x"24",x"18",x"00",x"00",x"42", -- 0x15E0
		x"42",x"42",x"42",x"5A",x"24",x"00",x"00",x"42", -- 0x15E8
		x"24",x"18",x"18",x"24",x"42",x"00",x"00",x"82", -- 0x15F0
		x"44",x"28",x"10",x"10",x"10",x"00",x"00",x"7E", -- 0x15F8
		x"04",x"08",x"10",x"20",x"7E",x"00",x"00",x"0E", -- 0x1600
		x"08",x"08",x"08",x"08",x"0E",x"00",x"00",x"00", -- 0x1608
		x"40",x"20",x"10",x"08",x"04",x"00",x"00",x"70", -- 0x1610
		x"10",x"10",x"10",x"10",x"70",x"00",x"00",x"10", -- 0x1618
		x"38",x"54",x"10",x"10",x"10",x"00",x"00",x"00", -- 0x1620
		x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"1C", -- 0x1628
		x"22",x"78",x"20",x"20",x"7E",x"00",x"00",x"00", -- 0x1630
		x"38",x"04",x"3C",x"44",x"3C",x"00",x"00",x"20", -- 0x1638
		x"20",x"3C",x"22",x"22",x"3C",x"00",x"00",x"00", -- 0x1640
		x"1C",x"20",x"20",x"20",x"1C",x"00",x"00",x"04", -- 0x1648
		x"04",x"3C",x"44",x"44",x"3C",x"00",x"00",x"00", -- 0x1650
		x"38",x"44",x"78",x"40",x"3C",x"00",x"00",x"0C", -- 0x1658
		x"10",x"18",x"10",x"10",x"10",x"00",x"00",x"00", -- 0x1660
		x"3C",x"44",x"44",x"3C",x"04",x"38",x"00",x"40", -- 0x1668
		x"40",x"78",x"44",x"44",x"44",x"00",x"00",x"10", -- 0x1670
		x"00",x"30",x"10",x"10",x"38",x"00",x"00",x"04", -- 0x1678
		x"00",x"04",x"04",x"04",x"24",x"18",x"00",x"20", -- 0x1680
		x"28",x"30",x"30",x"28",x"24",x"00",x"00",x"10", -- 0x1688
		x"10",x"10",x"10",x"10",x"0C",x"00",x"00",x"00", -- 0x1690
		x"68",x"54",x"54",x"54",x"54",x"00",x"00",x"00", -- 0x1698
		x"78",x"44",x"44",x"44",x"44",x"00",x"00",x"00", -- 0x16A0
		x"38",x"44",x"44",x"44",x"38",x"00",x"00",x"00", -- 0x16A8
		x"78",x"44",x"44",x"78",x"40",x"40",x"00",x"00", -- 0x16B0
		x"3C",x"44",x"44",x"3C",x"04",x"06",x"00",x"00", -- 0x16B8
		x"1C",x"20",x"20",x"20",x"20",x"00",x"00",x"00", -- 0x16C0
		x"38",x"40",x"38",x"04",x"78",x"00",x"00",x"10", -- 0x16C8
		x"38",x"10",x"10",x"10",x"0C",x"00",x"00",x"00", -- 0x16D0
		x"44",x"44",x"44",x"44",x"38",x"00",x"00",x"00", -- 0x16D8
		x"44",x"44",x"28",x"28",x"10",x"00",x"00",x"00", -- 0x16E0
		x"44",x"54",x"54",x"54",x"28",x"00",x"00",x"00", -- 0x16E8
		x"44",x"28",x"10",x"28",x"44",x"00",x"00",x"00", -- 0x16F0
		x"44",x"44",x"44",x"3C",x"04",x"38",x"00",x"00", -- 0x16F8
		x"7C",x"08",x"10",x"20",x"7C",x"00",x"00",x"0E", -- 0x1700
		x"08",x"30",x"08",x"08",x"0E",x"00",x"00",x"08", -- 0x1708
		x"08",x"08",x"08",x"08",x"08",x"00",x"00",x"70", -- 0x1710
		x"10",x"0C",x"10",x"10",x"70",x"00",x"00",x"14", -- 0x1718
		x"28",x"00",x"00",x"00",x"00",x"00",x"3C",x"42", -- 0x1720
		x"99",x"A1",x"A1",x"99",x"42",x"3C",x"00",x"C0", -- 0x1728
		x"02",x"2C",x"00",x"00",x"00",x"F7",x"FD",x"21", -- 0x1730
		x"02",x"00",x"FD",x"39",x"FD",x"7E",x"00",x"D3", -- 0x1738
		x"99",x"FD",x"7E",x"01",x"E6",x"3F",x"5F",x"16", -- 0x1740
		x"00",x"21",x"04",x"00",x"39",x"7E",x"E6",x"01", -- 0x1748
		x"0F",x"0F",x"E6",x"C0",x"4F",x"06",x"00",x"7B", -- 0x1750
		x"B1",x"67",x"7A",x"B0",x"7C",x"D3",x"99",x"C9", -- 0x1758
		x"3E",x"01",x"F5",x"33",x"21",x"05",x"00",x"39", -- 0x1760
		x"4E",x"23",x"46",x"C5",x"CD",x"36",x"17",x"F1", -- 0x1768
		x"33",x"11",x"00",x"00",x"21",x"06",x"00",x"39", -- 0x1770
		x"7B",x"96",x"7A",x"23",x"9E",x"D0",x"21",x"02", -- 0x1778
		x"00",x"39",x"7E",x"23",x"66",x"6F",x"19",x"7E", -- 0x1780
		x"D3",x"98",x"26",x"0A",x"7C",x"C6",x"FF",x"67", -- 0x1788
		x"B7",x"20",x"F9",x"13",x"18",x"DE",x"21",x"24", -- 0x1790
		x"44",x"34",x"3E",x"1F",x"FD",x"21",x"24",x"44", -- 0x1798
		x"FD",x"96",x"00",x"D0",x"21",x"24",x"44",x"36", -- 0x17A0
		x"00",x"21",x"25",x"44",x"34",x"3E",x"17",x"FD", -- 0x17A8
		x"21",x"25",x"44",x"FD",x"96",x"00",x"D0",x"21", -- 0x17B0
		x"25",x"44",x"36",x"17",x"C9",x"1E",x"00",x"21", -- 0x17B8
		x"2E",x"17",x"16",x"00",x"19",x"66",x"D5",x"E5", -- 0x17C0
		x"33",x"7B",x"F5",x"33",x"CD",x"1A",x"14",x"F1", -- 0x17C8
		x"D1",x"1C",x"7B",x"D6",x"08",x"38",x"E8",x"3E", -- 0x17D0
		x"01",x"F5",x"33",x"21",x"00",x"00",x"E5",x"CD", -- 0x17D8
		x"36",x"17",x"F1",x"33",x"11",x"00",x"00",x"3E", -- 0x17E0
		x"00",x"D3",x"98",x"13",x"7A",x"D6",x"01",x"38", -- 0x17E8
		x"F6",x"21",x"2E",x"14",x"01",x"00",x"03",x"C5", -- 0x17F0
		x"01",x"00",x"01",x"C5",x"E5",x"CD",x"60",x"17", -- 0x17F8
		x"F1",x"F1",x"26",x"01",x"E3",x"33",x"21",x"00", -- 0x1800
		x"04",x"E5",x"CD",x"36",x"17",x"F1",x"33",x"11", -- 0x1808
		x"00",x"00",x"3E",x"00",x"D3",x"98",x"13",x"7A", -- 0x1810
		x"D6",x"04",x"38",x"F6",x"21",x"25",x"44",x"36", -- 0x1818
		x"00",x"21",x"24",x"44",x"36",x"00",x"21",x"26", -- 0x1820
		x"44",x"36",x"0F",x"21",x"27",x"44",x"36",x"07", -- 0x1828
		x"3E",x"01",x"F5",x"33",x"21",x"00",x"08",x"E5", -- 0x1830
		x"CD",x"36",x"17",x"F1",x"33",x"11",x"00",x"00", -- 0x1838
		x"3E",x"20",x"D3",x"98",x"13",x"7A",x"D6",x"03", -- 0x1840
		x"38",x"F6",x"C9",x"3B",x"21",x"05",x"00",x"39", -- 0x1848
		x"7E",x"E6",x"0F",x"07",x"07",x"07",x"07",x"E6", -- 0x1850
		x"F0",x"67",x"FD",x"21",x"04",x"00",x"FD",x"39", -- 0x1858
		x"FD",x"7E",x"00",x"E6",x"0F",x"B4",x"33",x"F5", -- 0x1860
		x"33",x"FD",x"21",x"03",x"00",x"FD",x"39",x"FD", -- 0x1868
		x"7E",x"00",x"E6",x"0F",x"B4",x"57",x"1E",x"07", -- 0x1870
		x"D5",x"CD",x"1A",x"14",x"26",x"01",x"E3",x"33", -- 0x1878
		x"21",x"00",x"0B",x"E5",x"CD",x"36",x"17",x"F1", -- 0x1880
		x"33",x"16",x"00",x"21",x"00",x"00",x"39",x"7E", -- 0x1888
		x"D3",x"98",x"14",x"7A",x"D6",x"20",x"38",x"F3", -- 0x1890
		x"21",x"05",x"00",x"39",x"7E",x"32",x"26",x"44", -- 0x1898
		x"21",x"04",x"00",x"39",x"7E",x"32",x"27",x"44", -- 0x18A0
		x"33",x"C9",x"3E",x"01",x"F5",x"33",x"21",x"00", -- 0x18A8
		x"08",x"E5",x"CD",x"36",x"17",x"F1",x"33",x"11", -- 0x18B0
		x"00",x"00",x"3E",x"20",x"D3",x"98",x"13",x"7A", -- 0x18B8
		x"D6",x"03",x"38",x"F6",x"C9",x"21",x"02",x"00", -- 0x18C0
		x"39",x"7E",x"E6",x"1F",x"32",x"24",x"44",x"21", -- 0x18C8
		x"03",x"00",x"39",x"7E",x"32",x"25",x"44",x"3E", -- 0x18D0
		x"17",x"FD",x"21",x"25",x"44",x"FD",x"96",x"00", -- 0x18D8
		x"D0",x"21",x"25",x"44",x"36",x"17",x"C9",x"21", -- 0x18E0
		x"02",x"00",x"39",x"7E",x"E6",x"1F",x"32",x"24", -- 0x18E8
		x"44",x"21",x"03",x"00",x"39",x"7E",x"32",x"25", -- 0x18F0
		x"44",x"3E",x"17",x"FD",x"21",x"25",x"44",x"FD", -- 0x18F8
		x"96",x"00",x"30",x"05",x"21",x"25",x"44",x"36", -- 0x1900
		x"17",x"FD",x"21",x"25",x"44",x"FD",x"6E",x"00", -- 0x1908
		x"26",x"00",x"29",x"29",x"29",x"29",x"29",x"5D", -- 0x1910
		x"7C",x"C6",x"08",x"57",x"FD",x"21",x"24",x"44", -- 0x1918
		x"FD",x"6E",x"00",x"26",x"00",x"19",x"EB",x"3E", -- 0x1920
		x"01",x"F5",x"33",x"D5",x"CD",x"36",x"17",x"F1", -- 0x1928
		x"33",x"21",x"04",x"00",x"39",x"7E",x"D3",x"98", -- 0x1930
		x"C3",x"96",x"17",x"21",x"02",x"00",x"39",x"7E", -- 0x1938
		x"D6",x"0A",x"20",x"10",x"21",x"24",x"44",x"36", -- 0x1940
		x"00",x"3A",x"25",x"44",x"D6",x"17",x"D0",x"21", -- 0x1948
		x"25",x"44",x"34",x"C9",x"21",x"02",x"00",x"39", -- 0x1950
		x"7E",x"F5",x"33",x"3A",x"25",x"44",x"F5",x"33", -- 0x1958
		x"3A",x"24",x"44",x"F5",x"33",x"CD",x"E7",x"18", -- 0x1960
		x"F1",x"33",x"C9",x"21",x"24",x"44",x"5E",x"16", -- 0x1968
		x"00",x"21",x"00",x"0B",x"19",x"EB",x"21",x"03", -- 0x1970
		x"00",x"39",x"7E",x"E6",x"0F",x"07",x"07",x"07", -- 0x1978
		x"07",x"E6",x"F0",x"21",x"27",x"44",x"B6",x"47", -- 0x1980
		x"C5",x"3E",x"01",x"F5",x"33",x"D5",x"CD",x"36", -- 0x1988
		x"17",x"F1",x"33",x"C1",x"78",x"D3",x"98",x"21", -- 0x1990
		x"02",x"00",x"39",x"7E",x"F5",x"33",x"3A",x"25", -- 0x1998
		x"44",x"F5",x"33",x"3A",x"24",x"44",x"F5",x"33", -- 0x19A0
		x"CD",x"E7",x"18",x"F1",x"33",x"C9",x"C1",x"E1", -- 0x19A8
		x"E5",x"C5",x"56",x"E5",x"D5",x"33",x"CD",x"3B", -- 0x19B0
		x"19",x"33",x"E1",x"23",x"7E",x"B7",x"20",x"F2", -- 0x19B8
		x"C9",x"C1",x"E1",x"E5",x"C5",x"AF",x"47",x"4F", -- 0x19C0
		x"ED",x"B1",x"21",x"FF",x"FF",x"ED",x"42",x"C9", -- 0x19C8
		x"F1",x"E1",x"D1",x"D5",x"E5",x"F5",x"44",x"4D", -- 0x19D0
		x"AF",x"6F",x"B0",x"06",x"10",x"20",x"04",x"06", -- 0x19D8
		x"08",x"79",x"29",x"CB",x"11",x"17",x"30",x"01", -- 0x19E0
		x"19",x"10",x"F7",x"C9",x"DD",x"E5",x"DD",x"21", -- 0x19E8
		x"00",x"00",x"DD",x"39",x"21",x"FA",x"FF",x"39", -- 0x19F0
		x"F9",x"21",x"0A",x"00",x"39",x"4D",x"44",x"23", -- 0x19F8
		x"23",x"DD",x"75",x"FE",x"DD",x"74",x"FF",x"69", -- 0x1A00
		x"60",x"23",x"23",x"5E",x"23",x"56",x"21",x"0E", -- 0x1A08
		x"00",x"39",x"DD",x"75",x"FC",x"DD",x"74",x"FD", -- 0x1A10
		x"DD",x"6E",x"FC",x"DD",x"66",x"FD",x"7E",x"23", -- 0x1A18
		x"66",x"6F",x"C5",x"E5",x"D5",x"CD",x"D0",x"19", -- 0x1A20
		x"F1",x"F1",x"55",x"5C",x"C1",x"DD",x"6E",x"FE", -- 0x1A28
		x"DD",x"66",x"FF",x"72",x"23",x"73",x"69",x"60", -- 0x1A30
		x"23",x"23",x"DD",x"75",x"FE",x"DD",x"74",x"FF", -- 0x1A38
		x"69",x"60",x"23",x"23",x"7E",x"DD",x"77",x"FA", -- 0x1A40
		x"23",x"7E",x"DD",x"77",x"FB",x"D1",x"E1",x"E5", -- 0x1A48
		x"D5",x"23",x"23",x"5E",x"23",x"56",x"69",x"60", -- 0x1A50
		x"7E",x"23",x"66",x"6F",x"C5",x"E5",x"D5",x"CD", -- 0x1A58
		x"D0",x"19",x"F1",x"F1",x"C1",x"DD",x"7E",x"FA", -- 0x1A60
		x"85",x"57",x"DD",x"7E",x"FB",x"8C",x"5F",x"DD", -- 0x1A68
		x"6E",x"FE",x"DD",x"66",x"FF",x"72",x"23",x"73", -- 0x1A70
		x"69",x"60",x"23",x"23",x"E3",x"69",x"60",x"23", -- 0x1A78
		x"23",x"5E",x"23",x"56",x"69",x"60",x"23",x"7E", -- 0x1A80
		x"DD",x"77",x"FE",x"DD",x"6E",x"FC",x"DD",x"66", -- 0x1A88
		x"FD",x"23",x"66",x"D5",x"C5",x"DD",x"5E",x"FE", -- 0x1A90
		x"2E",x"00",x"55",x"06",x"08",x"29",x"30",x"01", -- 0x1A98
		x"19",x"10",x"FA",x"C1",x"D1",x"19",x"EB",x"E1", -- 0x1AA0
		x"E5",x"73",x"23",x"72",x"D1",x"E1",x"E5",x"D5", -- 0x1AA8
		x"5E",x"69",x"60",x"23",x"66",x"C5",x"2E",x"00", -- 0x1AB0
		x"55",x"06",x"08",x"29",x"30",x"01",x"19",x"10", -- 0x1AB8
		x"FA",x"C1",x"EB",x"DD",x"6E",x"FC",x"DD",x"66", -- 0x1AC0
		x"FD",x"23",x"E5",x"FD",x"E1",x"69",x"60",x"7E", -- 0x1AC8
		x"DD",x"77",x"FA",x"DD",x"6E",x"FC",x"DD",x"66", -- 0x1AD0
		x"FD",x"23",x"7E",x"D5",x"C5",x"5F",x"DD",x"66", -- 0x1AD8
		x"FA",x"2E",x"00",x"55",x"06",x"08",x"29",x"30", -- 0x1AE0
		x"01",x"19",x"10",x"FA",x"C1",x"D1",x"FD",x"75", -- 0x1AE8
		x"00",x"FD",x"74",x"01",x"DD",x"6E",x"FC",x"DD", -- 0x1AF0
		x"66",x"FD",x"23",x"23",x"23",x"E3",x"DD",x"6E", -- 0x1AF8
		x"FC",x"DD",x"66",x"FD",x"23",x"E5",x"FD",x"E1", -- 0x1B00
		x"DD",x"6E",x"FC",x"DD",x"66",x"FD",x"23",x"7E", -- 0x1B08
		x"23",x"66",x"6F",x"19",x"FD",x"75",x"00",x"FD", -- 0x1B10
		x"74",x"01",x"BF",x"ED",x"52",x"3E",x"00",x"17", -- 0x1B18
		x"E1",x"E5",x"77",x"59",x"50",x"0A",x"4F",x"DD", -- 0x1B20
		x"6E",x"FC",x"DD",x"66",x"FD",x"66",x"D5",x"59", -- 0x1B28
		x"2E",x"00",x"55",x"06",x"08",x"29",x"30",x"01", -- 0x1B30
		x"19",x"10",x"FA",x"D1",x"4D",x"44",x"79",x"12", -- 0x1B38
		x"13",x"78",x"12",x"C1",x"E1",x"E5",x"C5",x"36", -- 0x1B40
		x"00",x"DD",x"7E",x"04",x"DD",x"86",x"08",x"6F", -- 0x1B48
		x"DD",x"7E",x"05",x"DD",x"8E",x"09",x"67",x"DD", -- 0x1B50
		x"7E",x"06",x"DD",x"8E",x"0A",x"5F",x"DD",x"7E", -- 0x1B58
		x"07",x"DD",x"8E",x"0B",x"57",x"DD",x"F9",x"DD", -- 0x1B60
		x"E1",x"C9",x"5E",x"0A",x"6A",x"0A",x"76",x"0A", -- 0x1B68
		x"82",x"0A",x"8E",x"0A",x"9A",x"0A",x"A6",x"0A", -- 0x1B70
		x"B2",x"0A",x"01",x"10",x"00",x"78",x"B1",x"28", -- 0x1B78
		x"08",x"11",x"28",x"44",x"21",x"6A",x"1B",x"ED", -- 0x1B80
		x"B0",x"C9",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B88
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B90
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BA8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BB0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BD8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C08
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C10
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C28
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C30
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C38
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C40
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C48
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C80
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C88
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C90
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CA8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CB0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CD8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D08
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D10
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D28
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D30
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D38
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D40
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D48
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D80
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D88
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D90
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DA8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DB0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DD8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E08
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E10
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E28
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E30
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E38
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E40
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E48
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E80
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E88
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E90
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1EA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1EA8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1EB0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1EB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1EC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1EC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1ED0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1ED8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1EE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1EE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1EF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1EF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F08
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F10
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F28
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F30
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F38
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F40
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F48
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F80
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F88
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F90
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FA8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FB0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FD8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF"  -- 0x1FF8
	);

begin

	process(clk)
	begin
		if rising_edge(clk) then
			data <= ROM(to_integer(unsigned(addr)));
		end if;
	end process;
end RTL;
